module sigmoidFracData
(
	input	            clka,
	input		[7:0]	addra,
	input				ena,
	output		[13:0]	douta
);
reg [13:0] DATA;
assign	douta = DATA;
always@(posedge clka) begin
    if(ena) begin
        case(addra)
            8'd0 : DATA <= 14'd3128;
            8'd1 : DATA <= 14'd4292;
            8'd2 : DATA <= 14'd5889;
            8'd3 : DATA <= 14'd8081;
            8'd4 : DATA <= 14'd1109;
            8'd5 : DATA <= 14'd1522;
            8'd6 : DATA <= 14'd2088;
            8'd7 : DATA <= 14'd2865;
            8'd8 : DATA <= 14'd3931;
            8'd9 : DATA <= 14'd5395;
            8'd10 : DATA <= 14'd7403;
            8'd11 : DATA <= 14'd1016;
            8'd12 : DATA <= 14'd1394;
            8'd13 : DATA <= 14'd1913;
            8'd14 : DATA <= 14'd2624;
            8'd15 : DATA <= 14'd3601;
            8'd16 : DATA <= 14'd4942;
            8'd17 : DATA <= 14'd6781;
            8'd18 : DATA <= 14'd9305;
            8'd19 : DATA <= 14'd1277;
            8'd20 : DATA <= 14'd1752;
            8'd21 : DATA <= 14'd2404;
            8'd22 : DATA <= 14'd3299;
            8'd23 : DATA <= 14'd4527;
            8'd24 : DATA <= 14'd6211;
            8'd25 : DATA <= 14'd8523;
            8'd26 : DATA <= 14'd1170;
            8'd27 : DATA <= 14'd1605;
            8'd28 : DATA <= 14'd2202;
            8'd29 : DATA <= 14'd3022;
            8'd30 : DATA <= 14'd4147;
            8'd31 : DATA <= 14'd5690;
            8'd32 : DATA <= 14'd7807;
            8'd33 : DATA <= 14'd1071;
            8'd34 : DATA <= 14'd1470;
            8'd35 : DATA <= 14'd2017;
            8'd36 : DATA <= 14'd2768;
            8'd37 : DATA <= 14'd3798;
            8'd38 : DATA <= 14'd5212;
            8'd39 : DATA <= 14'd7152;
            8'd40 : DATA <= 14'd9814;
            8'd41 : DATA <= 14'd1347;
            8'd42 : DATA <= 14'd1848;
            8'd43 : DATA <= 14'd2536;
            8'd44 : DATA <= 14'd3479;
            8'd45 : DATA <= 14'd4774;
            8'd46 : DATA <= 14'd6551;
            8'd47 : DATA <= 14'd8990;
            8'd48 : DATA <= 14'd1234;
            8'd49 : DATA <= 14'd1693;
            8'd50 : DATA <= 14'd2323;
            8'd51 : DATA <= 14'd3187;
            8'd52 : DATA <= 14'd4373;
            8'd53 : DATA <= 14'd6001;
            8'd54 : DATA <= 14'd8235;
            8'd55 : DATA <= 14'd1130;
            8'd56 : DATA <= 14'd1550;
            8'd57 : DATA <= 14'd2128;
            8'd58 : DATA <= 14'd2919;
            8'd59 : DATA <= 14'd4006;
            8'd60 : DATA <= 14'd5497;
            8'd61 : DATA <= 14'd7543;
            8'd62 : DATA <= 14'd1035;
            8'd63 : DATA <= 14'd1420;
            8'd64 : DATA <= 14'd1949;
            8'd65 : DATA <= 14'd2674;
            8'd66 : DATA <= 14'd3668;
            8'd67 : DATA <= 14'd5033;
            8'd68 : DATA <= 14'd6905;
            8'd69 : DATA <= 14'd9472;
            8'd70 : DATA <= 14'd1299;
            8'd71 : DATA <= 14'd1782;
            8'd72 : DATA <= 14'd2444;
            8'd73 : DATA <= 14'd3350;
            8'd74 : DATA <= 14'd4591;
            8'd75 : DATA <= 14'd6290;
            8'd76 : DATA <= 14'd8610;
            8'd77 : DATA <= 14'd1178;
            8'd78 : DATA <= 14'd1609;
            8'd79 : DATA <= 14'd2195;
            8'd80 : DATA <= 14'd2987;
            8'd81 : DATA <= 14'd4054;
            8'd82 : DATA <= 14'd5480;
            8'd83 : DATA <= 14'd7369;
            8'd84 : DATA <= 14'd9842;
            8'd85 : DATA <= 14'd1303;
            8'd86 : DATA <= 14'd1705;
            8'd87 : DATA <= 14'd2200;
            8'd88 : DATA <= 14'd2790;
            8'd89 : DATA <= 14'd3469;
            8'd90 : DATA <= 14'd4216;
            8'd91 : DATA <= 14'd5000;
            8'd92 : DATA <= 14'd5784;
            8'd93 : DATA <= 14'd6531;
            8'd94 : DATA <= 14'd7210;
            8'd95 : DATA <= 14'd7800;
            8'd96 : DATA <= 14'd8295;
            8'd97 : DATA <= 14'd8697;
            8'd98 : DATA <= 14'd9016;
            8'd99 : DATA <= 14'd9263;
            8'd100 : DATA <= 14'd9452;
            8'd101 : DATA <= 14'd9595;
            8'd102 : DATA <= 14'd9701;
            8'd103 : DATA <= 14'd9781;
            8'd104 : DATA <= 14'd9839;
            8'd105 : DATA <= 14'd9882;
            8'd106 : DATA <= 14'd9914;
            8'd107 : DATA <= 14'd9937;
            8'd108 : DATA <= 14'd9954;
            8'd109 : DATA <= 14'd9966;
            8'd110 : DATA <= 14'd9976;
            8'd111 : DATA <= 14'd9982;
            8'd112 : DATA <= 14'd9987;
            8'd113 : DATA <= 14'd9991;
            8'd114 : DATA <= 14'd9993;
            8'd115 : DATA <= 14'd9995;
            8'd116 : DATA <= 14'd9996;
            8'd117 : DATA <= 14'd9997;
            8'd118 : DATA <= 14'd9998;
            8'd119 : DATA <= 14'd9999;
            8'd120 : DATA <= 14'd9999;
            8'd121 : DATA <= 14'd9999;
            8'd122 : DATA <= 14'd9999;
            8'd123 : DATA <= 14'd1000;
            8'd124 : DATA <= 14'd1000;
            8'd125 : DATA <= 14'd1000;
            8'd126 : DATA <= 14'd1000;
            8'd127 : DATA <= 14'd1000;
            8'd128 : DATA <= 14'd1000;
            8'd129 : DATA <= 14'd1000;
            8'd130 : DATA <= 14'd1000;
            8'd131 : DATA <= 14'd1000;
            8'd132 : DATA <= 14'd1000;
            8'd133 : DATA <= 14'd1000;
            8'd134 : DATA <= 14'd1000;
            8'd135 : DATA <= 14'd1000;
            8'd136 : DATA <= 14'd1000;
            8'd137 : DATA <= 14'd1000;
            8'd138 : DATA <= 14'd1000;
            8'd139 : DATA <= 14'd1000;
            8'd140 : DATA <= 14'd1000;
            8'd141 : DATA <= 14'd1000;
            8'd142 : DATA <= 14'd1000;
            8'd143 : DATA <= 14'd1000;
            8'd144 : DATA <= 14'd1000;
            8'd145 : DATA <= 14'd1000;
            8'd146 : DATA <= 14'd1000;
            8'd147 : DATA <= 14'd1000;
            8'd148 : DATA <= 14'd1000;
            8'd149 : DATA <= 14'd1000;
            8'd150 : DATA <= 14'd1000;
            8'd151 : DATA <= 14'd1000;
            8'd152 : DATA <= 14'd1000;
            8'd153 : DATA <= 14'd1000;
            8'd154 : DATA <= 14'd1000;
            8'd155 : DATA <= 14'd1000;
            8'd156 : DATA <= 14'd1000;
            8'd157 : DATA <= 14'd1000;
            8'd158 : DATA <= 14'd1000;
            8'd159 : DATA <= 14'd1000;
            8'd160 : DATA <= 14'd1000;
            8'd161 : DATA <= 14'd1000;
            8'd162 : DATA <= 14'd1000;
            8'd163 : DATA <= 14'd1000;
            8'd164 : DATA <= 14'd1000;
            8'd165 : DATA <= 14'd1000;
            8'd166 : DATA <= 14'd1000;
            8'd167 : DATA <= 14'd1000;
            8'd168 : DATA <= 14'd1000;
            8'd169 : DATA <= 14'd1000;
            8'd170 : DATA <= 14'd1000;
            8'd171 : DATA <= 14'd1000;
            8'd172 : DATA <= 14'd1000;
            8'd173 : DATA <= 14'd1000;
            8'd174 : DATA <= 14'd1000;
            8'd175 : DATA <= 14'd1000;
            8'd176 : DATA <= 14'd1000;
            8'd177 : DATA <= 14'd1000;
            8'd178 : DATA <= 14'd1000;
            8'd179 : DATA <= 14'd1000;
            8'd180 : DATA <= 14'd1000;
            8'd181 : DATA <= 14'd1000;
            8'd182 : DATA <= 14'd1000;
            8'd183 : DATA <= 14'd1000;
            8'd184 : DATA <= 14'd1000;
            8'd185 : DATA <= 14'd1000;
            8'd186 : DATA <= 14'd1000;
            8'd187 : DATA <= 14'd1000;
            8'd188 : DATA <= 14'd1000;
            8'd189 : DATA <= 14'd1000;
            8'd190 : DATA <= 14'd1000;
            8'd191 : DATA <= 14'd1000;
            8'd192 : DATA <= 14'd1000;
            8'd193 : DATA <= 14'd1000;
            8'd194 : DATA <= 14'd1000;
            8'd195 : DATA <= 14'd1000;
            8'd196 : DATA <= 14'd1000;
            8'd197 : DATA <= 14'd1000;
            8'd198 : DATA <= 14'd1000;
            8'd199 : DATA <= 14'd1000;
            8'd200 : DATA <= 14'd1000;
            8'd201 : DATA <= 14'd1000;
            8'd202 : DATA <= 14'd1000;
            8'd203 : DATA <= 14'd1000;
            8'd204 : DATA <= 14'd1000;
            8'd205 : DATA <= 14'd1000;
            8'd206 : DATA <= 14'd1000;
            8'd207 : DATA <= 14'd1000;
            8'd208 : DATA <= 14'd1000;
            8'd209 : DATA <= 14'd1000;
            8'd210 : DATA <= 14'd1000;
            8'd211 : DATA <= 14'd1000;
            8'd212 : DATA <= 14'd1000;
            8'd213 : DATA <= 14'd1000;
            8'd214 : DATA <= 14'd1000;
            8'd215 : DATA <= 14'd1000;
            8'd216 : DATA <= 14'd1000;
            8'd217 : DATA <= 14'd1000;
            8'd218 : DATA <= 14'd1000;
            8'd219 : DATA <= 14'd1000;
            8'd220 : DATA <= 14'd1000;
            8'd221 : DATA <= 14'd1000;
            8'd222 : DATA <= 14'd1000;
            8'd223 : DATA <= 14'd1000;
            8'd224 : DATA <= 14'd1000;
            8'd225 : DATA <= 14'd1000;
            8'd226 : DATA <= 14'd1000;
            8'd227 : DATA <= 14'd1000;
            8'd228 : DATA <= 14'd1000;
            8'd229 : DATA <= 14'd1000;
            8'd230 : DATA <= 14'd1000;
            8'd231 : DATA <= 14'd1000;
            8'd232 : DATA <= 14'd1000;
            8'd233 : DATA <= 14'd1000;
            8'd234 : DATA <= 14'd1000;
            8'd235 : DATA <= 14'd1000;
            8'd236 : DATA <= 14'd1000;
            8'd237 : DATA <= 14'd1000;
            8'd238 : DATA <= 14'd1000;
            8'd239 : DATA <= 14'd1000;
            8'd240 : DATA <= 14'd1000;
            8'd241 : DATA <= 14'd1000;
            8'd242 : DATA <= 14'd1000;
            8'd243 : DATA <= 14'd1000;
            8'd244 : DATA <= 14'd1000;
            8'd245 : DATA <= 14'd1000;
            8'd246 : DATA <= 14'd1000;
            8'd247 : DATA <= 14'd1000;
            8'd248 : DATA <= 14'd1000;
            8'd249 : DATA <= 14'd1000;
            8'd250 : DATA <= 14'd1000;
            8'd251 : DATA <= 14'd1000;
            8'd252 : DATA <= 14'd1000;
            8'd253 : DATA <= 14'd1000;
            8'd254 : DATA <= 14'd1000;
            8'd255 : DATA <= 14'd1000;
            default:   DATA<= 0;
        endcase
    end
end
endmodule
