`timescale 1ns / 1ps

module uart_tx_path(
	input clk_i,
	input [7:0] uart_tx_data_i,	//待发送数据
	input uart_tx_en_i,			//发送发送使能信号
	output uart_tx_o,
	output uart_busy
);

parameter [13:0] BAUD_DIV     = 14'd433;//波特率时钟，115200bps，50Mhz/115200 - 1'b1=433
//波特率发生器，实际就是分配器
reg bps_start_en = 1'b0;
reg [13:0] baud_div = 14'd0;

assign uart_busy = bps_start_en;

always@(posedge clk_i)begin
    if(bps_start_en && baud_div < BAUD_DIV)	
        baud_div <= baud_div + 1'b1;
    else 
        baud_div <= 14'd0;
end

reg [9:0] uart_tx_data_r = 10'h3ff;
wire bps_en = (baud_div == BAUD_DIV);
reg [3:0] tx_cnt = 4'd0;
assign uart_tx_o = uart_tx_data_r[0];
always@(posedge clk_i)begin
//首先当发送使能有效，寄存数据
    if(uart_tx_en_i) begin
        bps_start_en <= 1'b1;
        tx_cnt <= 4'd0;
        uart_tx_data_r <= {1'b1,uart_tx_data_i[7:0],1'b0};
    end
    else if(!bps_start_en)begin//当bps_start_en为0让状态机处于停止状态
        uart_tx_data_r <= 10'h3ff;
        tx_cnt <= 4'd0;
    end
// 通过移位发送数据
    if(bps_en && tx_cnt < 4'd9)begin
         uart_tx_data_r <= {uart_tx_data_r[0],uart_tx_data_r[9:1]};
         tx_cnt <= tx_cnt + 1'b1;
    end
    else if(bps_en)begin
         bps_start_en <= 1'd0;
    end
end   

endmodule

