module Accel_Conv
#(
	parameter FM_ADDR_BIT=12,
	parameter WEIGHT_AXI_ADDR_BIT=14,
	parameter WEIGHTBUF_ADDR_BIT=7,
	parameter BIASBUF_ADDR_BIT=7,
	
	parameter FM_DEPTH=4096,
	parameter WEIGHTBUF_DEPTH=128,
	parameter BIASBUF_DEPTH=128,
	
	parameter LINEBUFFER_LEN1=15,
	parameter LINEBUFFER_LEN2=13,
	parameter LINEBUFFER_LEN3=26,
	parameter LINEBUFFER_LEN4=52,
	parameter LINEBUFFER_LEN5=104,
	parameter LINEBUFFER_LEN6=208,

	parameter C_S_AXI_DATA_WIDTH = 32,
	parameter C_S_AXI_ADDR_WIDTH = 7,
	
	parameter IFM_RAM_STYLE="block",
	parameter WEIGHT_RAM_STYLE="distributed",
	parameter BIAS_RAM_STYLE="distributed",
	parameter OFM_RAM_STYLE="block"
)
(
	input clk,
	input rst,
    output yolo_layer_finish,  
	output resize_load,
	input  yolo_clr,
	// output [31:0] pwm0_reg,
	// output [31:0] pwm1_reg,
	input e203_clk,
	input e203_rst_n,
	input [5:0]  send_addr,
	output [31:0] send_data,
	
	// axi-lite interface
	
	//dma_read interface
	output	[31:0]	dma_raddr,
	output			dma_rareq,
	output	[15:0]	dma_rsize,
	input 			dma_rbusy,
	input	[63:0]  dma_rdata,
	input 			dma_rvalid,
	output			dma_rready,

	//dma_write interface
	output [31:0]   dma_waddr,
	output 			dma_wareq,
	output [15:0]	dma_wsize,
	input  			dma_wbusy,
	output [63:0]   dma_wdata,
	input  			dma_wvalid,
	output 			dma_wready
);
	wire ap_done;
	wire yolo_layer_en;

	//accel control reg
	wire [31:0] reg_0;
	wire [31:0] reg_1;
	wire [31:0] reg_2;
	wire [31:0] reg_3;
	//dma control reg
	wire [31:0] reg_4;
	wire [31:0] reg_5;
	wire [31:0] reg_6;
	wire [31:0] reg_7;

	wire [31:0]	dma_slave_addr;
	wire [15:0]	dma_slave_len;
	wire [31:0]	dma_master_addr;
	wire [15:0] dma_master_len;
	assign dma_slave_addr = reg_4;
	assign dma_slave_len  = {reg_5[18:3]};
	assign dma_master_addr = reg_6;
	assign dma_master_len = {reg_7[18:3]};


	// reg 0
	wire			recv_enable;
	wire			send_enable;
	wire			conv_start;
	wire			pool_enable;
	wire			first_conv;
	wire			last_conv;
	wire			ifmbuf_sel;
	wire			task_valid;
	wire	[1:0]	axis_buf_sel;
	wire	[2:0]	sel;
	wire	[1:0]	ofm_send_sel;
	wire			pool_stride_sel;
	wire	[7:0]	row;
	wire			relu_type_sel;
	
	// reg 1 reg 2
	wire	[15:0]	scale;
    wire	[3:0]	shift;
	wire	[7:0]	zero_point_in;
	wire	[7:0]	zero_point_out;
	wire	[7:0]	zero_point_act;
	
	// reg 2 reg 3
	wire	[WEIGHTBUF_ADDR_BIT-1:0]	weightbuf_read_addr_in;
	wire	[BIASBUF_ADDR_BIT-1:0]		biasbuf_read_addr_in;
	
	// reg 0
	assign recv_enable     =reg_0[0];
	assign send_enable     =reg_0[1];
	assign axis_buf_sel    =reg_0[3:2];
	assign conv_start      =reg_0[4];
	assign pool_enable     =reg_0[5];
	assign first_conv      =reg_0[6];
	assign last_conv       =reg_0[7];
	assign ifmbuf_sel      =reg_0[8];
	assign task_valid      =reg_0[9];
	assign sel             =reg_0[12:10];
	assign ofm_send_sel    =reg_0[14:13];
	assign pool_stride_sel =reg_0[15];
	assign relu_type_sel   =reg_0[16];
	assign row             =reg_0[31:24];

	// reg 1 reg 2
	assign scale          =reg_1[15:0];
	assign shift          =reg_1[19:16];
	assign zero_point_in  =reg_2[7:0];
	assign zero_point_out =reg_2[15:8];
	assign zero_point_act =reg_2[23:16];
	
	// reg 3
	assign weightbuf_read_addr_in =reg_3[WEIGHTBUF_ADDR_BIT-1:0];
	assign biasbuf_read_addr_in   =reg_3[16+BIASBUF_ADDR_BIT-1:16];

	// global parameter
	wire	[8:0]				conv_row;
	wire	[8:0]				conv_col;
	wire	[8:0]				pool_row;
	wire	[8:0]				pool_col;
	wire	[FM_ADDR_BIT-1:0]	conv_addr_len;
	wire	[FM_ADDR_BIT-1:0]	pool_addr_len;
	wire	[FM_ADDR_BIT-1:0]	ofm_addr_start;
	wire	[FM_ADDR_BIT-1:0]	ofm_addr_end;

	// ifm buffer
	wire	[FM_ADDR_BIT+1-2:0]	ifmbuf_bram_addr_write;
	wire	[FM_ADDR_BIT+1-2:0]	ifmbuf_bram_addr_read;
	wire ifmbuf_bram_en_write;
	
	// weight buffer
	wire								weightbuf_waddr_clear;
	wire								weightbuf_bram_en_write;
	wire	[WEIGHTBUF_ADDR_BIT-1:0]	weightbuf_read_addr;
	assign weightbuf_read_addr=weightbuf_read_addr_in;
	
	// bias buffer
	wire							biasbuf_waddr_clear;
	wire							biasbuf_bram_en_write;
	wire	[BIASBUF_ADDR_BIT-1:0]	biasbuf_read_addr;
	assign biasbuf_read_addr=biasbuf_read_addr_in;
	
	// ofm buffer
	wire						ofmbuf_bram_en_write;
	wire	[FM_ADDR_BIT-1:0]	ofmbuf_bram_write_addr;
	wire	[FM_ADDR_BIT-1:0]	ofmbuf_bram_read_addr;
	wire	[FM_ADDR_BIT-1:0]	ofm_after_quant_addr;
	wire						ofm_after_quant_valid;
	wire						ofm_after_quant_done;
	wire	[FM_ADDR_BIT-1:0]	ofm_after_pool_addr;
	wire						ofm_after_pool_valid;
	wire						ofm_after_pool_zero;
	wire						ofm_after_pool_done;
	assign ofmbuf_bram_en_write=(pool_enable==1'b1)?ofm_after_pool_valid:ofm_after_quant_valid;
	assign ofmbuf_bram_write_addr=(pool_enable==1'b1)?ofm_after_pool_addr:ofm_after_quant_addr;
	
	// acc
	wire						acc_read_en;
	wire						acc_write_en;
	wire	[FM_ADDR_BIT-1:0]	acc_read_addr;
	wire	[FM_ADDR_BIT-1:0]	acc_write_addr;
	wire						acc_prev_data_zero;
	wire						acc_curr_data_zero;
	assign acc_prev_data_zero=first_conv;
	
	// pool
	wire pool_zero_out;
	assign pool_zero_out=ofm_after_pool_zero;
	
	// ifm data port
	wire [7:0] ifm_in_0;
	wire [7:0] ifm_in_1;
	wire [7:0] ifm_in_2;
	wire [7:0] ifm_in_3;
	wire [7:0] ifm_in_4;
	wire [7:0] ifm_in_5;
	wire [7:0] ifm_in_6;
	wire [7:0] ifm_in_7;
	
	// weight data port
	wire [7:0] weight_in_0;
	wire [7:0] weight_in_1;
	wire [7:0] weight_in_2;
	wire [7:0] weight_in_3;
	wire [7:0] weight_in_4;
	wire [7:0] weight_in_5;
	wire [7:0] weight_in_6;
	wire [7:0] weight_in_7;
	
	// bias data port
	wire [17:0] bias_in;
	
	// ofm bundle
	wire [63:0] ofm_out_bundle;
	
	// control signal
	wire			recv_done;
	wire			send_done;
	wire			recv_running;
	wire			send_running;
	wire			write_enable;
	wire	[15:0]	write_addr;
	wire	[63:0]	write_data;
	wire	[15:0]	read_addr;
	wire	[63:0]	read_data;
	
	wire	conv_shutdown;
	wire	conv_done_t;
	reg		conv_done;
	assign conv_done_t=(pool_enable==1'b1)?ofm_after_pool_done:ofm_after_quant_done;
	always@(posedge clk) begin
		conv_done<=conv_done_t;
	end
	assign weightbuf_waddr_clear=task_valid;
	assign biasbuf_waddr_clear=task_valid;
	
	// interface
	wire	[15:0]		write_addr_ifm;
	wire	[63:0]		write_data_ifm;
	wire				write_enable_ifm;
	wire	[15:0]		write_addr_weight;
	wire	[63:0]		write_data_weight;
	wire				write_enable_weight;
	wire	[15:0]		write_addr_bias;
	wire	[63:0]		write_data_bias;
	wire				write_enable_bias;
	wire	[15:0]		write_addr_leakyrelu;
	wire	[63:0]		write_data_leakyrelu;
	wire				write_enable_leakyrelu;

	assign ifmbuf_bram_addr_write  =write_addr_ifm[FM_ADDR_BIT+1-2:0];
	assign ifmbuf_bram_en_write    =write_enable_ifm;
	assign ifm_in_0                =write_data_ifm[7:0];
	assign ifm_in_1                =write_data_ifm[15:8];
	assign ifm_in_2                =write_data_ifm[23:16];
	assign ifm_in_3                =write_data_ifm[31:24];
	assign ifm_in_4                =write_data_ifm[39:32];
	assign ifm_in_5                =write_data_ifm[47:40];
	assign ifm_in_6                =write_data_ifm[55:48];
	assign ifm_in_7                =write_data_ifm[63:56];

	assign weightbuf_bram_en_write =write_enable_weight;
	assign weight_in_0             =write_data_weight[7:0];
	assign weight_in_1             =write_data_weight[15:8];
	assign weight_in_2             =write_data_weight[23:16];
	assign weight_in_3             =write_data_weight[31:24];
	assign weight_in_4             =write_data_weight[39:32];
	assign weight_in_5             =write_data_weight[47:40];
	assign weight_in_6             =write_data_weight[55:48];
	assign weight_in_7             =write_data_weight[63:56];

	assign biasbuf_bram_en_write   =write_enable_bias;
	assign bias_in                 =write_data_bias;
	
	assign ofmbuf_bram_read_addr   =read_addr[FM_ADDR_BIT-1:0];
	assign read_data               =ofm_out_bundle;

	global_para_gen
	#(
		.FM_ADDR_BIT(FM_ADDR_BIT),
		.LINEBUFFER_LEN1(LINEBUFFER_LEN1),
		.LINEBUFFER_LEN2(LINEBUFFER_LEN2),
		.LINEBUFFER_LEN3(LINEBUFFER_LEN3),
		.LINEBUFFER_LEN4(LINEBUFFER_LEN4),
		.LINEBUFFER_LEN5(LINEBUFFER_LEN5),
		.LINEBUFFER_LEN6(LINEBUFFER_LEN6)
	)
	u_global_para_gen
	(
		.clk(clk),
		.sel(sel),
		.row(row),
		.ofm_send_sel(ofm_send_sel),
		.pool_enable((~pool_stride_sel)&&pool_enable),
		
		.conv_row(conv_row),
		.conv_col(conv_col),
		.pool_row(pool_row),
		.pool_col(pool_col),
		
		.conv_addr_len(conv_addr_len),
		.pool_addr_len(pool_addr_len),
		.ofm_addr_start(ofm_addr_start),
		.ofm_addr_end(ofm_addr_end)
	);

	// wire [3:0]  conv_layer_cnt;
    // wire [31:0] delay_cnt;
    // wire conv_layer_finish;
	yolov3_tiny_ctrl u_yolov3_tiny_ctrl(
		.clk                      ( clk             ),
		.rst                      ( rst             ),
		.yolo_layer_finish        (yolo_layer_finish),
		// .conv_layer_cnt           (conv_layer_cnt),
		// .delay_cnt                (delay_cnt),
		// .conv_layer_finish        (conv_layer_finish),
		.yolo_clr                 (yolo_clr         ),
		.ap_done                  ( ap_done         ),
		.yolo_en                  ( yolo_layer_en   ),
		.resize_load              ( resize_load     ),
		.reg0                     ( reg_0           ),
		.reg1                     ( reg_1           ),
		.reg2                     ( reg_2           ),
		.reg3                     ( reg_3           ),
		.reg4                     ( reg_4           ),
		.reg5                     ( reg_5           ),
		.reg6                     ( reg_6           ),
		.reg7                     ( reg_7           )
	);

	generate_ctrl_signal inst_generate_ctrl_signal (
		.clk           (clk),
		.rst           (rst),
		.recv_enable   (recv_enable),
		.send_enable   (send_enable),
		.conv_start    (conv_start),
		.recv_done     (recv_done),
		.send_done     (send_done),
		.conv_done     (conv_done),
		.recv_running  (recv_running),
		.send_running  (send_running),
		.conv_shutdown (conv_shutdown),
		.task_valid    (task_valid),
		.ap_done       (ap_done)
	);

	interface_dma_slave#(
		.ADDR_BIT ( 16 )
	)u_interface_dma_slave(
		.clk           ( clk         ),
		.rst_n         ( !rst       ),
		.recv_enable   ( recv_enable ),
		.recv_done     ( recv_done   ),
		.dma_addr      ( dma_slave_addr    ),
		.dma_len       ( dma_slave_len     ),
		.dma_raddr    ( dma_raddr  ),
		.dma_rareq    ( dma_rareq  ),
		.dma_rsize    ( dma_rsize  ),
		.dma_rbusy    ( dma_rbusy  ),
		.dma_rdata    ( dma_rdata  ),
		.dma_rvalid   ( dma_rvalid ),
		.dma_rready   ( dma_rready ),
		.write_addr    ( write_addr  ),
		.write_data    ( write_data  ),
		.write_enable  ( write_enable)
	);


	inferface_dma_master#(
		.ADDR_BIT    ( 16 )
	)u_inferface_dma_master(
		.clk         ( clk         ),
		.rst_n       ( !rst        ),
		.send_enable ( send_enable ),
		.send_done   ( send_done   ),
		.dma_addr    ( dma_master_addr    ),
		.dma_len     ( dma_master_len     ),
		.dma_waddr  ( dma_waddr  ),
		.dma_wareq  ( dma_wareq  ),
		.dma_wsize  ( dma_wsize  ),
		.dma_wbusy  ( dma_wbusy  ),
		.dma_wdata  ( dma_wdata  ),
		.dma_wvalid ( dma_wvalid ),
		.dma_wready ( dma_wready ),
		.addr_end    ( {{4'b0000},ofm_addr_end}    ),
		.addr_start  ( {{4'b0000},ofm_addr_start}  ),
		.read_addr   ( read_addr   ),
		.read_data   ( read_data   )
	);


	axis_buf_sel #(
		.DMA_ADDR_BIT(16)
	) inst_axis_buf_sel (
		.axis_buf_sel           (axis_buf_sel),
		.write_addr             (write_addr),
		.write_data             (write_data),
		.write_enable           (write_enable),

		.write_addr_ifm         (write_addr_ifm),
		.write_data_ifm         (write_data_ifm),
		.write_enable_ifm       (write_enable_ifm),

		.write_addr_weight      (write_addr_weight),
		.write_data_weight      (write_data_weight),
		.write_enable_weight    (write_enable_weight),

		.write_addr_bias        (write_addr_bias),
		.write_data_bias        (write_data_bias),
		.write_enable_bias      (write_enable_bias),

		.write_addr_leakyrelu   (write_addr_leakyrelu),
		.write_data_leakyrelu   (write_data_leakyrelu),
		.write_enable_leakyrelu (write_enable_leakyrelu)
	);

	global_data_beat
	#(.ADDR_BIT(FM_ADDR_BIT))
	u_global_data_beat
	(
		.clk(clk),
		.shutdown(conv_shutdown),
		
		.conv_addr_len(conv_addr_len),
		.pool_addr_len(pool_addr_len),
		.conv_col(conv_col),
		.conv_row(conv_row),
		.pool_stride_sel(pool_stride_sel),
		
		.ifmbuf_bram_addr_read(ifmbuf_bram_addr_read),
		
		.acc_read_en(acc_read_en),
		.acc_write_en(acc_write_en),
		.acc_read_addr(acc_read_addr),
		.acc_write_addr(acc_write_addr),
		.acc_curr_data_zero(acc_curr_data_zero),
		
		.ofm_after_quant_addr(ofm_after_quant_addr),
		.ofm_after_quant_valid(ofm_after_quant_valid),
		.ofm_after_quant_done(ofm_after_quant_done),
		
		.ofm_after_pool_addr(ofm_after_pool_addr),
		.ofm_after_pool_valid(ofm_after_pool_valid),
		.ofm_after_pool_zero(ofm_after_pool_zero),
		.ofm_after_pool_done(ofm_after_pool_done)
	);

	accel_top
	#(
		.IFMBUF_ADDR_BIT(FM_ADDR_BIT+1),
		.WEIGHTBUF_ADDR_BIT(WEIGHTBUF_ADDR_BIT),
		.BIASBUF_ADDR_BIT(BIASBUF_ADDR_BIT),
		.ACC_ADDR_BIT(FM_ADDR_BIT),
		.OFMBUF_ADDR_BIT(FM_ADDR_BIT),
		
		.IFMBUF_DEPTH(FM_DEPTH*2),
		.WEIGHTBUF_DEPTH(WEIGHTBUF_DEPTH),
		.BIASBUF_DEPTH(BIASBUF_DEPTH),
		.ACC_DEPTH(FM_DEPTH),
		.OFMBUF_DEPTH(FM_DEPTH),
		
		.LINEBUFFER_LEN1(LINEBUFFER_LEN1),
		.LINEBUFFER_LEN2(LINEBUFFER_LEN2),
		.LINEBUFFER_LEN3(LINEBUFFER_LEN3),
		.LINEBUFFER_LEN4(LINEBUFFER_LEN4),
		.LINEBUFFER_LEN5(LINEBUFFER_LEN5),
		.LINEBUFFER_LEN6(LINEBUFFER_LEN6),
		
		.IFM_RAM_STYLE(IFM_RAM_STYLE),
		.WEIGHT_RAM_STYLE(WEIGHT_RAM_STYLE),
		.BIAS_RAM_STYLE(BIAS_RAM_STYLE),
		.OFM_RAM_STYLE(OFM_RAM_STYLE)
	)
	u_accel_top
	(
		.clk(clk),
		.rst(rst),
		
		.sel(sel),
		.relu_type_sel(relu_type_sel),
		.pool_enable(pool_enable),
		
		.ifmbuf_bram_addr_write(ifmbuf_bram_addr_write),
		.ifmbuf_bram_addr_read(ifmbuf_bram_addr_read),
		.ifmbuf_bram_en_write(ifmbuf_bram_en_write),
		.ifmbuf_sel(ifmbuf_sel),
		
		.weightbuf_waddr_clear(weightbuf_waddr_clear),
		.weightbuf_bram_en_write(weightbuf_bram_en_write),
		.weightbuf_read_addr(weightbuf_read_addr),
		
		.biasbuf_waddr_clear(biasbuf_waddr_clear),
		.biasbuf_bram_en_write(biasbuf_bram_en_write),
		.biasbuf_read_addr(biasbuf_read_addr),
		
		.acc_read_en(acc_read_en),
		.acc_write_en(acc_write_en),
		.acc_read_addr(acc_read_addr),
		.acc_write_addr(acc_write_addr),
		.acc_prev_data_zero(acc_prev_data_zero),
		.acc_curr_data_zero(acc_curr_data_zero),
		
		.pool_zero_out(pool_zero_out),
		
		.ofmbuf_bram_en_write(ofmbuf_bram_en_write),
		.ofmbuf_bram_write_addr(ofmbuf_bram_write_addr),
		.ofmbuf_bram_read_addr(ofmbuf_bram_read_addr),
		
		.scale(scale),
		.shift(shift),
		.zero_point_in(zero_point_in),
		.zero_point_out(zero_point_out),
		.zero_point_act(zero_point_act),
		
		.ifm_in_0(ifm_in_0),
		.ifm_in_1(ifm_in_1),
		.ifm_in_2(ifm_in_2),
		.ifm_in_3(ifm_in_3),
		.ifm_in_4(ifm_in_4),
		.ifm_in_5(ifm_in_5),
		.ifm_in_6(ifm_in_6),
		.ifm_in_7(ifm_in_7),
		
		.weight_in_0(weight_in_0),
		.weight_in_1(weight_in_1),
		.weight_in_2(weight_in_2),
		.weight_in_3(weight_in_3),
		.weight_in_4(weight_in_4),
		.weight_in_5(weight_in_5),
		.weight_in_6(weight_in_6),
		.weight_in_7(weight_in_7),

		.write_addr_leakyrelu(write_addr_leakyrelu),
		.write_data_leakyrelu(write_data_leakyrelu),
		.write_enable_leakyrelu(write_enable_leakyrelu),
		
		.bias_in(bias_in),
		.bias_valid(last_conv),
		
		.ofm_out_bundle(ofm_out_bundle)
	);	

module_yolo_layer u_module_yolo_layer(
    .clk               ( clk               ),
    .rst               ( rst              ),
	.e203_clk          (e203_clk           ),
	.e203_rst_n        (e203_rst_n         ),
	.yolo_clr          ( yolo_clr          ),
    .dma_wdata        ( dma_wdata        ),
    .dma_wvalid       ( dma_wvalid       ),
    .dma_wbusy        ( dma_wbusy        ),
    .yolo_layer_en     ( yolo_layer_en     ),
    .yolo_layer_finish ( yolo_layer_finish ),
	.send_addr         (send_addr          ),
	.send_data         (send_data          )
);


endmodule