module sigmoidExpData
(
	input	            clka,
	input		[7:0]	addra,
	input				ena,
	output		[3:0]	douta
);
reg [3:0] DATA;
assign	douta = DATA;
always@(posedge clka) begin
    if(ena) begin
        case(addra)
            8'd0 : DATA <= 4'd13;
            8'd1 : DATA <= 4'd13;
            8'd2 : DATA <= 4'd13;
            8'd3 : DATA <= 4'd13;
            8'd4 : DATA <= 4'd12;
            8'd5 : DATA <= 4'd12;
            8'd6 : DATA <= 4'd12;
            8'd7 : DATA <= 4'd12;
            8'd8 : DATA <= 4'd12;
            8'd9 : DATA <= 4'd12;
            8'd10 : DATA <= 4'd12;
            8'd11 : DATA <= 4'd11;
            8'd12 : DATA <= 4'd11;
            8'd13 : DATA <= 4'd11;
            8'd14 : DATA <= 4'd11;
            8'd15 : DATA <= 4'd11;
            8'd16 : DATA <= 4'd11;
            8'd17 : DATA <= 4'd11;
            8'd18 : DATA <= 4'd11;
            8'd19 : DATA <= 4'd10;
            8'd20 : DATA <= 4'd10;
            8'd21 : DATA <= 4'd10;
            8'd22 : DATA <= 4'd10;
            8'd23 : DATA <= 4'd10;
            8'd24 : DATA <= 4'd10;
            8'd25 : DATA <= 4'd10;
            8'd26 : DATA <= 4'd9;
            8'd27 : DATA <= 4'd9;
            8'd28 : DATA <= 4'd9;
            8'd29 : DATA <= 4'd9;
            8'd30 : DATA <= 4'd9;
            8'd31 : DATA <= 4'd9;
            8'd32 : DATA <= 4'd9;
            8'd33 : DATA <= 4'd8;
            8'd34 : DATA <= 4'd8;
            8'd35 : DATA <= 4'd8;
            8'd36 : DATA <= 4'd8;
            8'd37 : DATA <= 4'd8;
            8'd38 : DATA <= 4'd8;
            8'd39 : DATA <= 4'd8;
            8'd40 : DATA <= 4'd8;
            8'd41 : DATA <= 4'd7;
            8'd42 : DATA <= 4'd7;
            8'd43 : DATA <= 4'd7;
            8'd44 : DATA <= 4'd7;
            8'd45 : DATA <= 4'd7;
            8'd46 : DATA <= 4'd7;
            8'd47 : DATA <= 4'd7;
            8'd48 : DATA <= 4'd6;
            8'd49 : DATA <= 4'd6;
            8'd50 : DATA <= 4'd6;
            8'd51 : DATA <= 4'd6;
            8'd52 : DATA <= 4'd6;
            8'd53 : DATA <= 4'd6;
            8'd54 : DATA <= 4'd6;
            8'd55 : DATA <= 4'd5;
            8'd56 : DATA <= 4'd5;
            8'd57 : DATA <= 4'd5;
            8'd58 : DATA <= 4'd5;
            8'd59 : DATA <= 4'd5;
            8'd60 : DATA <= 4'd5;
            8'd61 : DATA <= 4'd5;
            8'd62 : DATA <= 4'd4;
            8'd63 : DATA <= 4'd4;
            8'd64 : DATA <= 4'd4;
            8'd65 : DATA <= 4'd4;
            8'd66 : DATA <= 4'd4;
            8'd67 : DATA <= 4'd4;
            8'd68 : DATA <= 4'd4;
            8'd69 : DATA <= 4'd4;
            8'd70 : DATA <= 4'd3;
            8'd71 : DATA <= 4'd3;
            8'd72 : DATA <= 4'd3;
            8'd73 : DATA <= 4'd3;
            8'd74 : DATA <= 4'd3;
            8'd75 : DATA <= 4'd3;
            8'd76 : DATA <= 4'd3;
            8'd77 : DATA <= 4'd2;
            8'd78 : DATA <= 4'd2;
            8'd79 : DATA <= 4'd2;
            8'd80 : DATA <= 4'd2;
            8'd81 : DATA <= 4'd2;
            8'd82 : DATA <= 4'd2;
            8'd83 : DATA <= 4'd2;
            8'd84 : DATA <= 4'd2;
            8'd85 : DATA <= 4'd1;
            8'd86 : DATA <= 4'd1;
            8'd87 : DATA <= 4'd1;
            8'd88 : DATA <= 4'd1;
            8'd89 : DATA <= 4'd1;
            8'd90 : DATA <= 4'd1;
            8'd91 : DATA <= 4'd1;
            8'd92 : DATA <= 4'd1;
            8'd93 : DATA <= 4'd1;
            8'd94 : DATA <= 4'd1;
            8'd95 : DATA <= 4'd1;
            8'd96 : DATA <= 4'd1;
            8'd97 : DATA <= 4'd1;
            8'd98 : DATA <= 4'd1;
            8'd99 : DATA <= 4'd1;
            8'd100 : DATA <= 4'd1;
            8'd101 : DATA <= 4'd1;
            8'd102 : DATA <= 4'd1;
            8'd103 : DATA <= 4'd1;
            8'd104 : DATA <= 4'd1;
            8'd105 : DATA <= 4'd1;
            8'd106 : DATA <= 4'd1;
            8'd107 : DATA <= 4'd1;
            8'd108 : DATA <= 4'd1;
            8'd109 : DATA <= 4'd1;
            8'd110 : DATA <= 4'd1;
            8'd111 : DATA <= 4'd1;
            8'd112 : DATA <= 4'd1;
            8'd113 : DATA <= 4'd1;
            8'd114 : DATA <= 4'd1;
            8'd115 : DATA <= 4'd1;
            8'd116 : DATA <= 4'd1;
            8'd117 : DATA <= 4'd1;
            8'd118 : DATA <= 4'd1;
            8'd119 : DATA <= 4'd1;
            8'd120 : DATA <= 4'd1;
            8'd121 : DATA <= 4'd1;
            8'd122 : DATA <= 4'd1;
            8'd123 : DATA <= 4'd0;
            8'd124 : DATA <= 4'd0;
            8'd125 : DATA <= 4'd0;
            8'd126 : DATA <= 4'd0;
            8'd127 : DATA <= 4'd0;
            8'd128 : DATA <= 4'd0;
            8'd129 : DATA <= 4'd0;
            8'd130 : DATA <= 4'd0;
            8'd131 : DATA <= 4'd0;
            8'd132 : DATA <= 4'd0;
            8'd133 : DATA <= 4'd0;
            8'd134 : DATA <= 4'd0;
            8'd135 : DATA <= 4'd0;
            8'd136 : DATA <= 4'd0;
            8'd137 : DATA <= 4'd0;
            8'd138 : DATA <= 4'd0;
            8'd139 : DATA <= 4'd0;
            8'd140 : DATA <= 4'd0;
            8'd141 : DATA <= 4'd0;
            8'd142 : DATA <= 4'd0;
            8'd143 : DATA <= 4'd0;
            8'd144 : DATA <= 4'd0;
            8'd145 : DATA <= 4'd0;
            8'd146 : DATA <= 4'd0;
            8'd147 : DATA <= 4'd0;
            8'd148 : DATA <= 4'd0;
            8'd149 : DATA <= 4'd0;
            8'd150 : DATA <= 4'd0;
            8'd151 : DATA <= 4'd0;
            8'd152 : DATA <= 4'd0;
            8'd153 : DATA <= 4'd0;
            8'd154 : DATA <= 4'd0;
            8'd155 : DATA <= 4'd0;
            8'd156 : DATA <= 4'd0;
            8'd157 : DATA <= 4'd0;
            8'd158 : DATA <= 4'd0;
            8'd159 : DATA <= 4'd0;
            8'd160 : DATA <= 4'd0;
            8'd161 : DATA <= 4'd0;
            8'd162 : DATA <= 4'd0;
            8'd163 : DATA <= 4'd0;
            8'd164 : DATA <= 4'd0;
            8'd165 : DATA <= 4'd0;
            8'd166 : DATA <= 4'd0;
            8'd167 : DATA <= 4'd0;
            8'd168 : DATA <= 4'd0;
            8'd169 : DATA <= 4'd0;
            8'd170 : DATA <= 4'd0;
            8'd171 : DATA <= 4'd0;
            8'd172 : DATA <= 4'd0;
            8'd173 : DATA <= 4'd0;
            8'd174 : DATA <= 4'd0;
            8'd175 : DATA <= 4'd0;
            8'd176 : DATA <= 4'd0;
            8'd177 : DATA <= 4'd0;
            8'd178 : DATA <= 4'd0;
            8'd179 : DATA <= 4'd0;
            8'd180 : DATA <= 4'd0;
            8'd181 : DATA <= 4'd0;
            8'd182 : DATA <= 4'd0;
            8'd183 : DATA <= 4'd0;
            8'd184 : DATA <= 4'd0;
            8'd185 : DATA <= 4'd0;
            8'd186 : DATA <= 4'd0;
            8'd187 : DATA <= 4'd0;
            8'd188 : DATA <= 4'd0;
            8'd189 : DATA <= 4'd0;
            8'd190 : DATA <= 4'd0;
            8'd191 : DATA <= 4'd0;
            8'd192 : DATA <= 4'd0;
            8'd193 : DATA <= 4'd0;
            8'd194 : DATA <= 4'd0;
            8'd195 : DATA <= 4'd0;
            8'd196 : DATA <= 4'd0;
            8'd197 : DATA <= 4'd0;
            8'd198 : DATA <= 4'd0;
            8'd199 : DATA <= 4'd0;
            8'd200 : DATA <= 4'd0;
            8'd201 : DATA <= 4'd0;
            8'd202 : DATA <= 4'd0;
            8'd203 : DATA <= 4'd0;
            8'd204 : DATA <= 4'd0;
            8'd205 : DATA <= 4'd0;
            8'd206 : DATA <= 4'd0;
            8'd207 : DATA <= 4'd0;
            8'd208 : DATA <= 4'd0;
            8'd209 : DATA <= 4'd0;
            8'd210 : DATA <= 4'd0;
            8'd211 : DATA <= 4'd0;
            8'd212 : DATA <= 4'd0;
            8'd213 : DATA <= 4'd0;
            8'd214 : DATA <= 4'd0;
            8'd215 : DATA <= 4'd0;
            8'd216 : DATA <= 4'd0;
            8'd217 : DATA <= 4'd0;
            8'd218 : DATA <= 4'd0;
            8'd219 : DATA <= 4'd0;
            8'd220 : DATA <= 4'd0;
            8'd221 : DATA <= 4'd0;
            8'd222 : DATA <= 4'd0;
            8'd223 : DATA <= 4'd0;
            8'd224 : DATA <= 4'd0;
            8'd225 : DATA <= 4'd0;
            8'd226 : DATA <= 4'd0;
            8'd227 : DATA <= 4'd0;
            8'd228 : DATA <= 4'd0;
            8'd229 : DATA <= 4'd0;
            8'd230 : DATA <= 4'd0;
            8'd231 : DATA <= 4'd0;
            8'd232 : DATA <= 4'd0;
            8'd233 : DATA <= 4'd0;
            8'd234 : DATA <= 4'd0;
            8'd235 : DATA <= 4'd0;
            8'd236 : DATA <= 4'd0;
            8'd237 : DATA <= 4'd0;
            8'd238 : DATA <= 4'd0;
            8'd239 : DATA <= 4'd0;
            8'd240 : DATA <= 4'd0;
            8'd241 : DATA <= 4'd0;
            8'd242 : DATA <= 4'd0;
            8'd243 : DATA <= 4'd0;
            8'd244 : DATA <= 4'd0;
            8'd245 : DATA <= 4'd0;
            8'd246 : DATA <= 4'd0;
            8'd247 : DATA <= 4'd0;
            8'd248 : DATA <= 4'd0;
            8'd249 : DATA <= 4'd0;
            8'd250 : DATA <= 4'd0;
            8'd251 : DATA <= 4'd0;
            8'd252 : DATA <= 4'd0;
            8'd253 : DATA <= 4'd0;
            8'd254 : DATA <= 4'd0;
            8'd255 : DATA <= 4'd0;
            default:   DATA<= 0;
        endcase
    end
end
endmodule
