module CharOutput(
  input         clock,
  input         reset,
  input  [10:0] io_h_cnt,
  input  [10:0] io_v_cnt,
  input  [4:0]  io_class_voc_0,
  input  [4:0]  io_class_voc_1,
  input  [4:0]  io_class_voc_2,
  input  [4:0]  io_class_voc_3,
  input  [4:0]  io_class_voc_4,
  input  [10:0] io_rect_xleft_0,
  input  [10:0] io_rect_xleft_1,
  input  [10:0] io_rect_xleft_2,
  input  [10:0] io_rect_xleft_3,
  input  [10:0] io_rect_xleft_4,
  input  [10:0] io_rect_ytop_0,
  input  [10:0] io_rect_ytop_1,
  input  [10:0] io_rect_ytop_2,
  input  [10:0] io_rect_ytop_3,
  input  [10:0] io_rect_ytop_4,
  output        io_pixel,
  output        io_char_area_valid_0,
  output        io_char_area_valid_1,
  output        io_char_area_valid_2,
  output        io_char_area_valid_3,
  output        io_char_area_valid_4
);
  reg [11:0] dot_txt [0:4095]; // @[CharOutput.scala 105:20]
  wire  dot_txt_io_pixel_MPORT_en; // @[CharOutput.scala 105:20]
  wire [11:0] dot_txt_io_pixel_MPORT_addr; // @[CharOutput.scala 105:20]
  wire [11:0] dot_txt_io_pixel_MPORT_data; // @[CharOutput.scala 105:20]
  wire [6:0] _GEN_1 = 5'h1 == io_class_voc_0 ? 7'h3f : 7'h51; // @[CharOutput.scala 54:{24,24}]
  wire [6:0] _GEN_2 = 5'h2 == io_class_voc_0 ? 7'h24 : _GEN_1; // @[CharOutput.scala 54:{24,24}]
  wire [6:0] _GEN_3 = 5'h3 == io_class_voc_0 ? 7'h24 : _GEN_2; // @[CharOutput.scala 54:{24,24}]
  wire [6:0] _GEN_4 = 5'h4 == io_class_voc_0 ? 7'h36 : _GEN_3; // @[CharOutput.scala 54:{24,24}]
  wire [6:0] _GEN_5 = 5'h5 == io_class_voc_0 ? 7'h1b : _GEN_4; // @[CharOutput.scala 54:{24,24}]
  wire [6:0] _GEN_6 = 5'h6 == io_class_voc_0 ? 7'h1b : _GEN_5; // @[CharOutput.scala 54:{24,24}]
  wire [6:0] _GEN_7 = 5'h7 == io_class_voc_0 ? 7'h1b : _GEN_6; // @[CharOutput.scala 54:{24,24}]
  wire [6:0] _GEN_8 = 5'h8 == io_class_voc_0 ? 7'h2d : _GEN_7; // @[CharOutput.scala 54:{24,24}]
  wire [6:0] _GEN_9 = 5'h9 == io_class_voc_0 ? 7'h1b : _GEN_8; // @[CharOutput.scala 54:{24,24}]
  wire [6:0] _GEN_10 = 5'ha == io_class_voc_0 ? 7'h63 : _GEN_9; // @[CharOutput.scala 54:{24,24}]
  wire [6:0] _GEN_11 = 5'hb == io_class_voc_0 ? 7'h1b : _GEN_10; // @[CharOutput.scala 54:{24,24}]
  wire [6:0] _GEN_12 = 5'hc == io_class_voc_0 ? 7'h2d : _GEN_11; // @[CharOutput.scala 54:{24,24}]
  wire [6:0] _GEN_13 = 5'hd == io_class_voc_0 ? 7'h51 : _GEN_12; // @[CharOutput.scala 54:{24,24}]
  wire [6:0] _GEN_14 = 5'he == io_class_voc_0 ? 7'h36 : _GEN_13; // @[CharOutput.scala 54:{24,24}]
  wire [6:0] _GEN_15 = 5'hf == io_class_voc_0 ? 7'h63 : _GEN_14; // @[CharOutput.scala 54:{24,24}]
  wire [6:0] _GEN_16 = 5'h10 == io_class_voc_0 ? 7'h2d : _GEN_15; // @[CharOutput.scala 54:{24,24}]
  wire [6:0] _GEN_17 = 5'h11 == io_class_voc_0 ? 7'h24 : _GEN_16; // @[CharOutput.scala 54:{24,24}]
  wire [6:0] _GEN_18 = 5'h12 == io_class_voc_0 ? 7'h2d : _GEN_17; // @[CharOutput.scala 54:{24,24}]
  wire [6:0] char_area_width_0 = 5'h13 == io_class_voc_0 ? 7'h51 : _GEN_18; // @[CharOutput.scala 54:{24,24}]
  wire [10:0] _GEN_1618 = {{4'd0}, char_area_width_0}; // @[CharOutput.scala 57:45]
  wire [10:0] char_area_xright_0 = io_rect_xleft_0 + _GEN_1618; // @[CharOutput.scala 57:45]
  wire [10:0] char_area_ytop_0 = io_rect_ytop_0 - 11'h10; // @[CharOutput.scala 58:42]
  wire  in_area_h_0 = io_h_cnt < char_area_xright_0 & io_h_cnt >= io_rect_xleft_0; // @[CharOutput.scala 61:54]
  wire  in_area_v_0 = io_v_cnt >= char_area_ytop_0 & io_v_cnt < io_rect_ytop_0; // @[CharOutput.scala 62:53]
  wire  char_area_en_0 = in_area_h_0 & in_area_v_0; // @[CharOutput.scala 63:23]
  wire [6:0] _GEN_22 = 5'h1 == io_class_voc_1 ? 7'h3f : 7'h51; // @[CharOutput.scala 54:{24,24}]
  wire [6:0] _GEN_23 = 5'h2 == io_class_voc_1 ? 7'h24 : _GEN_22; // @[CharOutput.scala 54:{24,24}]
  wire [6:0] _GEN_24 = 5'h3 == io_class_voc_1 ? 7'h24 : _GEN_23; // @[CharOutput.scala 54:{24,24}]
  wire [6:0] _GEN_25 = 5'h4 == io_class_voc_1 ? 7'h36 : _GEN_24; // @[CharOutput.scala 54:{24,24}]
  wire [6:0] _GEN_26 = 5'h5 == io_class_voc_1 ? 7'h1b : _GEN_25; // @[CharOutput.scala 54:{24,24}]
  wire [6:0] _GEN_27 = 5'h6 == io_class_voc_1 ? 7'h1b : _GEN_26; // @[CharOutput.scala 54:{24,24}]
  wire [6:0] _GEN_28 = 5'h7 == io_class_voc_1 ? 7'h1b : _GEN_27; // @[CharOutput.scala 54:{24,24}]
  wire [6:0] _GEN_29 = 5'h8 == io_class_voc_1 ? 7'h2d : _GEN_28; // @[CharOutput.scala 54:{24,24}]
  wire [6:0] _GEN_30 = 5'h9 == io_class_voc_1 ? 7'h1b : _GEN_29; // @[CharOutput.scala 54:{24,24}]
  wire [6:0] _GEN_31 = 5'ha == io_class_voc_1 ? 7'h63 : _GEN_30; // @[CharOutput.scala 54:{24,24}]
  wire [6:0] _GEN_32 = 5'hb == io_class_voc_1 ? 7'h1b : _GEN_31; // @[CharOutput.scala 54:{24,24}]
  wire [6:0] _GEN_33 = 5'hc == io_class_voc_1 ? 7'h2d : _GEN_32; // @[CharOutput.scala 54:{24,24}]
  wire [6:0] _GEN_34 = 5'hd == io_class_voc_1 ? 7'h51 : _GEN_33; // @[CharOutput.scala 54:{24,24}]
  wire [6:0] _GEN_35 = 5'he == io_class_voc_1 ? 7'h36 : _GEN_34; // @[CharOutput.scala 54:{24,24}]
  wire [6:0] _GEN_36 = 5'hf == io_class_voc_1 ? 7'h63 : _GEN_35; // @[CharOutput.scala 54:{24,24}]
  wire [6:0] _GEN_37 = 5'h10 == io_class_voc_1 ? 7'h2d : _GEN_36; // @[CharOutput.scala 54:{24,24}]
  wire [6:0] _GEN_38 = 5'h11 == io_class_voc_1 ? 7'h24 : _GEN_37; // @[CharOutput.scala 54:{24,24}]
  wire [6:0] _GEN_39 = 5'h12 == io_class_voc_1 ? 7'h2d : _GEN_38; // @[CharOutput.scala 54:{24,24}]
  wire [6:0] char_area_width_1 = 5'h13 == io_class_voc_1 ? 7'h51 : _GEN_39; // @[CharOutput.scala 54:{24,24}]
  wire [10:0] _GEN_1619 = {{4'd0}, char_area_width_1}; // @[CharOutput.scala 57:45]
  wire [10:0] char_area_xright_1 = io_rect_xleft_1 + _GEN_1619; // @[CharOutput.scala 57:45]
  wire [10:0] char_area_ytop_1 = io_rect_ytop_1 - 11'h10; // @[CharOutput.scala 58:42]
  wire  in_area_h_1 = io_h_cnt < char_area_xright_1 & io_h_cnt >= io_rect_xleft_1; // @[CharOutput.scala 61:54]
  wire  in_area_v_1 = io_v_cnt >= char_area_ytop_1 & io_v_cnt < io_rect_ytop_1; // @[CharOutput.scala 62:53]
  wire  char_area_en_1 = in_area_h_1 & in_area_v_1; // @[CharOutput.scala 63:23]
  wire [6:0] _GEN_43 = 5'h1 == io_class_voc_2 ? 7'h3f : 7'h51; // @[CharOutput.scala 54:{24,24}]
  wire [6:0] _GEN_44 = 5'h2 == io_class_voc_2 ? 7'h24 : _GEN_43; // @[CharOutput.scala 54:{24,24}]
  wire [6:0] _GEN_45 = 5'h3 == io_class_voc_2 ? 7'h24 : _GEN_44; // @[CharOutput.scala 54:{24,24}]
  wire [6:0] _GEN_46 = 5'h4 == io_class_voc_2 ? 7'h36 : _GEN_45; // @[CharOutput.scala 54:{24,24}]
  wire [6:0] _GEN_47 = 5'h5 == io_class_voc_2 ? 7'h1b : _GEN_46; // @[CharOutput.scala 54:{24,24}]
  wire [6:0] _GEN_48 = 5'h6 == io_class_voc_2 ? 7'h1b : _GEN_47; // @[CharOutput.scala 54:{24,24}]
  wire [6:0] _GEN_49 = 5'h7 == io_class_voc_2 ? 7'h1b : _GEN_48; // @[CharOutput.scala 54:{24,24}]
  wire [6:0] _GEN_50 = 5'h8 == io_class_voc_2 ? 7'h2d : _GEN_49; // @[CharOutput.scala 54:{24,24}]
  wire [6:0] _GEN_51 = 5'h9 == io_class_voc_2 ? 7'h1b : _GEN_50; // @[CharOutput.scala 54:{24,24}]
  wire [6:0] _GEN_52 = 5'ha == io_class_voc_2 ? 7'h63 : _GEN_51; // @[CharOutput.scala 54:{24,24}]
  wire [6:0] _GEN_53 = 5'hb == io_class_voc_2 ? 7'h1b : _GEN_52; // @[CharOutput.scala 54:{24,24}]
  wire [6:0] _GEN_54 = 5'hc == io_class_voc_2 ? 7'h2d : _GEN_53; // @[CharOutput.scala 54:{24,24}]
  wire [6:0] _GEN_55 = 5'hd == io_class_voc_2 ? 7'h51 : _GEN_54; // @[CharOutput.scala 54:{24,24}]
  wire [6:0] _GEN_56 = 5'he == io_class_voc_2 ? 7'h36 : _GEN_55; // @[CharOutput.scala 54:{24,24}]
  wire [6:0] _GEN_57 = 5'hf == io_class_voc_2 ? 7'h63 : _GEN_56; // @[CharOutput.scala 54:{24,24}]
  wire [6:0] _GEN_58 = 5'h10 == io_class_voc_2 ? 7'h2d : _GEN_57; // @[CharOutput.scala 54:{24,24}]
  wire [6:0] _GEN_59 = 5'h11 == io_class_voc_2 ? 7'h24 : _GEN_58; // @[CharOutput.scala 54:{24,24}]
  wire [6:0] _GEN_60 = 5'h12 == io_class_voc_2 ? 7'h2d : _GEN_59; // @[CharOutput.scala 54:{24,24}]
  wire [6:0] char_area_width_2 = 5'h13 == io_class_voc_2 ? 7'h51 : _GEN_60; // @[CharOutput.scala 54:{24,24}]
  wire [10:0] _GEN_1620 = {{4'd0}, char_area_width_2}; // @[CharOutput.scala 57:45]
  wire [10:0] char_area_xright_2 = io_rect_xleft_2 + _GEN_1620; // @[CharOutput.scala 57:45]
  wire [10:0] char_area_ytop_2 = io_rect_ytop_2 - 11'h10; // @[CharOutput.scala 58:42]
  wire  in_area_h_2 = io_h_cnt < char_area_xright_2 & io_h_cnt >= io_rect_xleft_2; // @[CharOutput.scala 61:54]
  wire  in_area_v_2 = io_v_cnt >= char_area_ytop_2 & io_v_cnt < io_rect_ytop_2; // @[CharOutput.scala 62:53]
  wire  char_area_en_2 = in_area_h_2 & in_area_v_2; // @[CharOutput.scala 63:23]
  wire [6:0] _GEN_64 = 5'h1 == io_class_voc_3 ? 7'h3f : 7'h51; // @[CharOutput.scala 54:{24,24}]
  wire [6:0] _GEN_65 = 5'h2 == io_class_voc_3 ? 7'h24 : _GEN_64; // @[CharOutput.scala 54:{24,24}]
  wire [6:0] _GEN_66 = 5'h3 == io_class_voc_3 ? 7'h24 : _GEN_65; // @[CharOutput.scala 54:{24,24}]
  wire [6:0] _GEN_67 = 5'h4 == io_class_voc_3 ? 7'h36 : _GEN_66; // @[CharOutput.scala 54:{24,24}]
  wire [6:0] _GEN_68 = 5'h5 == io_class_voc_3 ? 7'h1b : _GEN_67; // @[CharOutput.scala 54:{24,24}]
  wire [6:0] _GEN_69 = 5'h6 == io_class_voc_3 ? 7'h1b : _GEN_68; // @[CharOutput.scala 54:{24,24}]
  wire [6:0] _GEN_70 = 5'h7 == io_class_voc_3 ? 7'h1b : _GEN_69; // @[CharOutput.scala 54:{24,24}]
  wire [6:0] _GEN_71 = 5'h8 == io_class_voc_3 ? 7'h2d : _GEN_70; // @[CharOutput.scala 54:{24,24}]
  wire [6:0] _GEN_72 = 5'h9 == io_class_voc_3 ? 7'h1b : _GEN_71; // @[CharOutput.scala 54:{24,24}]
  wire [6:0] _GEN_73 = 5'ha == io_class_voc_3 ? 7'h63 : _GEN_72; // @[CharOutput.scala 54:{24,24}]
  wire [6:0] _GEN_74 = 5'hb == io_class_voc_3 ? 7'h1b : _GEN_73; // @[CharOutput.scala 54:{24,24}]
  wire [6:0] _GEN_75 = 5'hc == io_class_voc_3 ? 7'h2d : _GEN_74; // @[CharOutput.scala 54:{24,24}]
  wire [6:0] _GEN_76 = 5'hd == io_class_voc_3 ? 7'h51 : _GEN_75; // @[CharOutput.scala 54:{24,24}]
  wire [6:0] _GEN_77 = 5'he == io_class_voc_3 ? 7'h36 : _GEN_76; // @[CharOutput.scala 54:{24,24}]
  wire [6:0] _GEN_78 = 5'hf == io_class_voc_3 ? 7'h63 : _GEN_77; // @[CharOutput.scala 54:{24,24}]
  wire [6:0] _GEN_79 = 5'h10 == io_class_voc_3 ? 7'h2d : _GEN_78; // @[CharOutput.scala 54:{24,24}]
  wire [6:0] _GEN_80 = 5'h11 == io_class_voc_3 ? 7'h24 : _GEN_79; // @[CharOutput.scala 54:{24,24}]
  wire [6:0] _GEN_81 = 5'h12 == io_class_voc_3 ? 7'h2d : _GEN_80; // @[CharOutput.scala 54:{24,24}]
  wire [6:0] char_area_width_3 = 5'h13 == io_class_voc_3 ? 7'h51 : _GEN_81; // @[CharOutput.scala 54:{24,24}]
  wire [10:0] _GEN_1621 = {{4'd0}, char_area_width_3}; // @[CharOutput.scala 57:45]
  wire [10:0] char_area_xright_3 = io_rect_xleft_3 + _GEN_1621; // @[CharOutput.scala 57:45]
  wire [10:0] char_area_ytop_3 = io_rect_ytop_3 - 11'h10; // @[CharOutput.scala 58:42]
  wire  in_area_h_3 = io_h_cnt < char_area_xright_3 & io_h_cnt >= io_rect_xleft_3; // @[CharOutput.scala 61:54]
  wire  in_area_v_3 = io_v_cnt >= char_area_ytop_3 & io_v_cnt < io_rect_ytop_3; // @[CharOutput.scala 62:53]
  wire  char_area_en_3 = in_area_h_3 & in_area_v_3; // @[CharOutput.scala 63:23]
  wire [6:0] _GEN_85 = 5'h1 == io_class_voc_4 ? 7'h3f : 7'h51; // @[CharOutput.scala 54:{24,24}]
  wire [6:0] _GEN_86 = 5'h2 == io_class_voc_4 ? 7'h24 : _GEN_85; // @[CharOutput.scala 54:{24,24}]
  wire [6:0] _GEN_87 = 5'h3 == io_class_voc_4 ? 7'h24 : _GEN_86; // @[CharOutput.scala 54:{24,24}]
  wire [6:0] _GEN_88 = 5'h4 == io_class_voc_4 ? 7'h36 : _GEN_87; // @[CharOutput.scala 54:{24,24}]
  wire [6:0] _GEN_89 = 5'h5 == io_class_voc_4 ? 7'h1b : _GEN_88; // @[CharOutput.scala 54:{24,24}]
  wire [6:0] _GEN_90 = 5'h6 == io_class_voc_4 ? 7'h1b : _GEN_89; // @[CharOutput.scala 54:{24,24}]
  wire [6:0] _GEN_91 = 5'h7 == io_class_voc_4 ? 7'h1b : _GEN_90; // @[CharOutput.scala 54:{24,24}]
  wire [6:0] _GEN_92 = 5'h8 == io_class_voc_4 ? 7'h2d : _GEN_91; // @[CharOutput.scala 54:{24,24}]
  wire [6:0] _GEN_93 = 5'h9 == io_class_voc_4 ? 7'h1b : _GEN_92; // @[CharOutput.scala 54:{24,24}]
  wire [6:0] _GEN_94 = 5'ha == io_class_voc_4 ? 7'h63 : _GEN_93; // @[CharOutput.scala 54:{24,24}]
  wire [6:0] _GEN_95 = 5'hb == io_class_voc_4 ? 7'h1b : _GEN_94; // @[CharOutput.scala 54:{24,24}]
  wire [6:0] _GEN_96 = 5'hc == io_class_voc_4 ? 7'h2d : _GEN_95; // @[CharOutput.scala 54:{24,24}]
  wire [6:0] _GEN_97 = 5'hd == io_class_voc_4 ? 7'h51 : _GEN_96; // @[CharOutput.scala 54:{24,24}]
  wire [6:0] _GEN_98 = 5'he == io_class_voc_4 ? 7'h36 : _GEN_97; // @[CharOutput.scala 54:{24,24}]
  wire [6:0] _GEN_99 = 5'hf == io_class_voc_4 ? 7'h63 : _GEN_98; // @[CharOutput.scala 54:{24,24}]
  wire [6:0] _GEN_100 = 5'h10 == io_class_voc_4 ? 7'h2d : _GEN_99; // @[CharOutput.scala 54:{24,24}]
  wire [6:0] _GEN_101 = 5'h11 == io_class_voc_4 ? 7'h24 : _GEN_100; // @[CharOutput.scala 54:{24,24}]
  wire [6:0] _GEN_102 = 5'h12 == io_class_voc_4 ? 7'h2d : _GEN_101; // @[CharOutput.scala 54:{24,24}]
  wire [6:0] char_area_width_4 = 5'h13 == io_class_voc_4 ? 7'h51 : _GEN_102; // @[CharOutput.scala 54:{24,24}]
  wire [10:0] _GEN_1622 = {{4'd0}, char_area_width_4}; // @[CharOutput.scala 57:45]
  wire [10:0] char_area_xright_4 = io_rect_xleft_4 + _GEN_1622; // @[CharOutput.scala 57:45]
  wire [10:0] char_area_ytop_4 = io_rect_ytop_4 - 11'h10; // @[CharOutput.scala 58:42]
  wire  in_area_h_4 = io_h_cnt < char_area_xright_4 & io_h_cnt >= io_rect_xleft_4; // @[CharOutput.scala 61:54]
  wire  in_area_v_4 = io_v_cnt >= char_area_ytop_4 & io_v_cnt < io_rect_ytop_4; // @[CharOutput.scala 62:53]
  wire  char_area_en_4 = in_area_h_4 & in_area_v_4; // @[CharOutput.scala 63:23]
  wire [5:0] _enc_T_1 = char_area_en_4 ? 6'h10 : 6'h20; // @[Mux.scala 47:70]
  wire [5:0] _enc_T_2 = char_area_en_3 ? 6'h8 : _enc_T_1; // @[Mux.scala 47:70]
  wire [5:0] _enc_T_3 = char_area_en_2 ? 6'h4 : _enc_T_2; // @[Mux.scala 47:70]
  wire [5:0] _enc_T_4 = char_area_en_1 ? 6'h2 : _enc_T_3; // @[Mux.scala 47:70]
  wire [5:0] enc = char_area_en_0 ? 6'h1 : _enc_T_4; // @[Mux.scala 47:70]
  wire  char_area_valid_5 = enc[5]; // @[OneHot.scala 82:30]
  wire [10:0] _char_index_0_T_1 = io_h_cnt - io_rect_xleft_0; // @[CharOutput.scala 82:48]
  wire [3:0] _GEN_114 = 7'h9 == _char_index_0_T_1[6:0] ? 4'h1 : 4'h0; // @[CharOutput.scala 82:{21,21}]
  wire [3:0] _GEN_115 = 7'ha == _char_index_0_T_1[6:0] ? 4'h1 : _GEN_114; // @[CharOutput.scala 82:{21,21}]
  wire [3:0] _GEN_116 = 7'hb == _char_index_0_T_1[6:0] ? 4'h1 : _GEN_115; // @[CharOutput.scala 82:{21,21}]
  wire [3:0] _GEN_117 = 7'hc == _char_index_0_T_1[6:0] ? 4'h1 : _GEN_116; // @[CharOutput.scala 82:{21,21}]
  wire [3:0] _GEN_118 = 7'hd == _char_index_0_T_1[6:0] ? 4'h1 : _GEN_117; // @[CharOutput.scala 82:{21,21}]
  wire [3:0] _GEN_119 = 7'he == _char_index_0_T_1[6:0] ? 4'h1 : _GEN_118; // @[CharOutput.scala 82:{21,21}]
  wire [3:0] _GEN_120 = 7'hf == _char_index_0_T_1[6:0] ? 4'h1 : _GEN_119; // @[CharOutput.scala 82:{21,21}]
  wire [3:0] _GEN_121 = 7'h10 == _char_index_0_T_1[6:0] ? 4'h1 : _GEN_120; // @[CharOutput.scala 82:{21,21}]
  wire [3:0] _GEN_122 = 7'h11 == _char_index_0_T_1[6:0] ? 4'h1 : _GEN_121; // @[CharOutput.scala 82:{21,21}]
  wire [3:0] _GEN_123 = 7'h12 == _char_index_0_T_1[6:0] ? 4'h2 : _GEN_122; // @[CharOutput.scala 82:{21,21}]
  wire [3:0] _GEN_124 = 7'h13 == _char_index_0_T_1[6:0] ? 4'h2 : _GEN_123; // @[CharOutput.scala 82:{21,21}]
  wire [3:0] _GEN_125 = 7'h14 == _char_index_0_T_1[6:0] ? 4'h2 : _GEN_124; // @[CharOutput.scala 82:{21,21}]
  wire [3:0] _GEN_126 = 7'h15 == _char_index_0_T_1[6:0] ? 4'h2 : _GEN_125; // @[CharOutput.scala 82:{21,21}]
  wire [3:0] _GEN_127 = 7'h16 == _char_index_0_T_1[6:0] ? 4'h2 : _GEN_126; // @[CharOutput.scala 82:{21,21}]
  wire [3:0] _GEN_128 = 7'h17 == _char_index_0_T_1[6:0] ? 4'h2 : _GEN_127; // @[CharOutput.scala 82:{21,21}]
  wire [3:0] _GEN_129 = 7'h18 == _char_index_0_T_1[6:0] ? 4'h2 : _GEN_128; // @[CharOutput.scala 82:{21,21}]
  wire [3:0] _GEN_130 = 7'h19 == _char_index_0_T_1[6:0] ? 4'h2 : _GEN_129; // @[CharOutput.scala 82:{21,21}]
  wire [3:0] _GEN_131 = 7'h1a == _char_index_0_T_1[6:0] ? 4'h2 : _GEN_130; // @[CharOutput.scala 82:{21,21}]
  wire [3:0] _GEN_132 = 7'h1b == _char_index_0_T_1[6:0] ? 4'h3 : _GEN_131; // @[CharOutput.scala 82:{21,21}]
  wire [3:0] _GEN_133 = 7'h1c == _char_index_0_T_1[6:0] ? 4'h3 : _GEN_132; // @[CharOutput.scala 82:{21,21}]
  wire [3:0] _GEN_134 = 7'h1d == _char_index_0_T_1[6:0] ? 4'h3 : _GEN_133; // @[CharOutput.scala 82:{21,21}]
  wire [3:0] _GEN_135 = 7'h1e == _char_index_0_T_1[6:0] ? 4'h3 : _GEN_134; // @[CharOutput.scala 82:{21,21}]
  wire [3:0] _GEN_136 = 7'h1f == _char_index_0_T_1[6:0] ? 4'h3 : _GEN_135; // @[CharOutput.scala 82:{21,21}]
  wire [3:0] _GEN_137 = 7'h20 == _char_index_0_T_1[6:0] ? 4'h3 : _GEN_136; // @[CharOutput.scala 82:{21,21}]
  wire [3:0] _GEN_138 = 7'h21 == _char_index_0_T_1[6:0] ? 4'h3 : _GEN_137; // @[CharOutput.scala 82:{21,21}]
  wire [3:0] _GEN_139 = 7'h22 == _char_index_0_T_1[6:0] ? 4'h3 : _GEN_138; // @[CharOutput.scala 82:{21,21}]
  wire [3:0] _GEN_140 = 7'h23 == _char_index_0_T_1[6:0] ? 4'h3 : _GEN_139; // @[CharOutput.scala 82:{21,21}]
  wire [3:0] _GEN_141 = 7'h24 == _char_index_0_T_1[6:0] ? 4'h4 : _GEN_140; // @[CharOutput.scala 82:{21,21}]
  wire [3:0] _GEN_142 = 7'h25 == _char_index_0_T_1[6:0] ? 4'h4 : _GEN_141; // @[CharOutput.scala 82:{21,21}]
  wire [3:0] _GEN_143 = 7'h26 == _char_index_0_T_1[6:0] ? 4'h4 : _GEN_142; // @[CharOutput.scala 82:{21,21}]
  wire [3:0] _GEN_144 = 7'h27 == _char_index_0_T_1[6:0] ? 4'h4 : _GEN_143; // @[CharOutput.scala 82:{21,21}]
  wire [3:0] _GEN_145 = 7'h28 == _char_index_0_T_1[6:0] ? 4'h4 : _GEN_144; // @[CharOutput.scala 82:{21,21}]
  wire [3:0] _GEN_146 = 7'h29 == _char_index_0_T_1[6:0] ? 4'h4 : _GEN_145; // @[CharOutput.scala 82:{21,21}]
  wire [3:0] _GEN_147 = 7'h2a == _char_index_0_T_1[6:0] ? 4'h4 : _GEN_146; // @[CharOutput.scala 82:{21,21}]
  wire [3:0] _GEN_148 = 7'h2b == _char_index_0_T_1[6:0] ? 4'h4 : _GEN_147; // @[CharOutput.scala 82:{21,21}]
  wire [3:0] _GEN_149 = 7'h2c == _char_index_0_T_1[6:0] ? 4'h4 : _GEN_148; // @[CharOutput.scala 82:{21,21}]
  wire [3:0] _GEN_150 = 7'h2d == _char_index_0_T_1[6:0] ? 4'h5 : _GEN_149; // @[CharOutput.scala 82:{21,21}]
  wire [3:0] _GEN_151 = 7'h2e == _char_index_0_T_1[6:0] ? 4'h5 : _GEN_150; // @[CharOutput.scala 82:{21,21}]
  wire [3:0] _GEN_152 = 7'h2f == _char_index_0_T_1[6:0] ? 4'h5 : _GEN_151; // @[CharOutput.scala 82:{21,21}]
  wire [3:0] _GEN_153 = 7'h30 == _char_index_0_T_1[6:0] ? 4'h5 : _GEN_152; // @[CharOutput.scala 82:{21,21}]
  wire [3:0] _GEN_154 = 7'h31 == _char_index_0_T_1[6:0] ? 4'h5 : _GEN_153; // @[CharOutput.scala 82:{21,21}]
  wire [3:0] _GEN_155 = 7'h32 == _char_index_0_T_1[6:0] ? 4'h5 : _GEN_154; // @[CharOutput.scala 82:{21,21}]
  wire [3:0] _GEN_156 = 7'h33 == _char_index_0_T_1[6:0] ? 4'h5 : _GEN_155; // @[CharOutput.scala 82:{21,21}]
  wire [3:0] _GEN_157 = 7'h34 == _char_index_0_T_1[6:0] ? 4'h5 : _GEN_156; // @[CharOutput.scala 82:{21,21}]
  wire [3:0] _GEN_158 = 7'h35 == _char_index_0_T_1[6:0] ? 4'h5 : _GEN_157; // @[CharOutput.scala 82:{21,21}]
  wire [3:0] _GEN_159 = 7'h36 == _char_index_0_T_1[6:0] ? 4'h6 : _GEN_158; // @[CharOutput.scala 82:{21,21}]
  wire [3:0] _GEN_160 = 7'h37 == _char_index_0_T_1[6:0] ? 4'h6 : _GEN_159; // @[CharOutput.scala 82:{21,21}]
  wire [3:0] _GEN_161 = 7'h38 == _char_index_0_T_1[6:0] ? 4'h6 : _GEN_160; // @[CharOutput.scala 82:{21,21}]
  wire [3:0] _GEN_162 = 7'h39 == _char_index_0_T_1[6:0] ? 4'h6 : _GEN_161; // @[CharOutput.scala 82:{21,21}]
  wire [3:0] _GEN_163 = 7'h3a == _char_index_0_T_1[6:0] ? 4'h6 : _GEN_162; // @[CharOutput.scala 82:{21,21}]
  wire [3:0] _GEN_164 = 7'h3b == _char_index_0_T_1[6:0] ? 4'h6 : _GEN_163; // @[CharOutput.scala 82:{21,21}]
  wire [3:0] _GEN_165 = 7'h3c == _char_index_0_T_1[6:0] ? 4'h6 : _GEN_164; // @[CharOutput.scala 82:{21,21}]
  wire [3:0] _GEN_166 = 7'h3d == _char_index_0_T_1[6:0] ? 4'h6 : _GEN_165; // @[CharOutput.scala 82:{21,21}]
  wire [3:0] _GEN_167 = 7'h3e == _char_index_0_T_1[6:0] ? 4'h6 : _GEN_166; // @[CharOutput.scala 82:{21,21}]
  wire [3:0] _GEN_168 = 7'h3f == _char_index_0_T_1[6:0] ? 4'h7 : _GEN_167; // @[CharOutput.scala 82:{21,21}]
  wire [3:0] _GEN_169 = 7'h40 == _char_index_0_T_1[6:0] ? 4'h7 : _GEN_168; // @[CharOutput.scala 82:{21,21}]
  wire [3:0] _GEN_170 = 7'h41 == _char_index_0_T_1[6:0] ? 4'h7 : _GEN_169; // @[CharOutput.scala 82:{21,21}]
  wire [3:0] _GEN_171 = 7'h42 == _char_index_0_T_1[6:0] ? 4'h7 : _GEN_170; // @[CharOutput.scala 82:{21,21}]
  wire [3:0] _GEN_172 = 7'h43 == _char_index_0_T_1[6:0] ? 4'h7 : _GEN_171; // @[CharOutput.scala 82:{21,21}]
  wire [3:0] _GEN_173 = 7'h44 == _char_index_0_T_1[6:0] ? 4'h7 : _GEN_172; // @[CharOutput.scala 82:{21,21}]
  wire [3:0] _GEN_174 = 7'h45 == _char_index_0_T_1[6:0] ? 4'h7 : _GEN_173; // @[CharOutput.scala 82:{21,21}]
  wire [3:0] _GEN_175 = 7'h46 == _char_index_0_T_1[6:0] ? 4'h7 : _GEN_174; // @[CharOutput.scala 82:{21,21}]
  wire [3:0] _GEN_176 = 7'h47 == _char_index_0_T_1[6:0] ? 4'h7 : _GEN_175; // @[CharOutput.scala 82:{21,21}]
  wire [3:0] _GEN_177 = 7'h48 == _char_index_0_T_1[6:0] ? 4'h8 : _GEN_176; // @[CharOutput.scala 82:{21,21}]
  wire [3:0] _GEN_178 = 7'h49 == _char_index_0_T_1[6:0] ? 4'h8 : _GEN_177; // @[CharOutput.scala 82:{21,21}]
  wire [3:0] _GEN_179 = 7'h4a == _char_index_0_T_1[6:0] ? 4'h8 : _GEN_178; // @[CharOutput.scala 82:{21,21}]
  wire [3:0] _GEN_180 = 7'h4b == _char_index_0_T_1[6:0] ? 4'h8 : _GEN_179; // @[CharOutput.scala 82:{21,21}]
  wire [3:0] _GEN_181 = 7'h4c == _char_index_0_T_1[6:0] ? 4'h8 : _GEN_180; // @[CharOutput.scala 82:{21,21}]
  wire [3:0] _GEN_182 = 7'h4d == _char_index_0_T_1[6:0] ? 4'h8 : _GEN_181; // @[CharOutput.scala 82:{21,21}]
  wire [3:0] _GEN_183 = 7'h4e == _char_index_0_T_1[6:0] ? 4'h8 : _GEN_182; // @[CharOutput.scala 82:{21,21}]
  wire [3:0] _GEN_184 = 7'h4f == _char_index_0_T_1[6:0] ? 4'h8 : _GEN_183; // @[CharOutput.scala 82:{21,21}]
  wire [3:0] _GEN_185 = 7'h50 == _char_index_0_T_1[6:0] ? 4'h8 : _GEN_184; // @[CharOutput.scala 82:{21,21}]
  wire [3:0] _GEN_186 = 7'h51 == _char_index_0_T_1[6:0] ? 4'h9 : _GEN_185; // @[CharOutput.scala 82:{21,21}]
  wire [3:0] _GEN_187 = 7'h52 == _char_index_0_T_1[6:0] ? 4'h9 : _GEN_186; // @[CharOutput.scala 82:{21,21}]
  wire [3:0] _GEN_188 = 7'h53 == _char_index_0_T_1[6:0] ? 4'h9 : _GEN_187; // @[CharOutput.scala 82:{21,21}]
  wire [3:0] _GEN_189 = 7'h54 == _char_index_0_T_1[6:0] ? 4'h9 : _GEN_188; // @[CharOutput.scala 82:{21,21}]
  wire [3:0] _GEN_190 = 7'h55 == _char_index_0_T_1[6:0] ? 4'h9 : _GEN_189; // @[CharOutput.scala 82:{21,21}]
  wire [3:0] _GEN_191 = 7'h56 == _char_index_0_T_1[6:0] ? 4'h9 : _GEN_190; // @[CharOutput.scala 82:{21,21}]
  wire [3:0] _GEN_192 = 7'h57 == _char_index_0_T_1[6:0] ? 4'h9 : _GEN_191; // @[CharOutput.scala 82:{21,21}]
  wire [3:0] _GEN_193 = 7'h58 == _char_index_0_T_1[6:0] ? 4'h9 : _GEN_192; // @[CharOutput.scala 82:{21,21}]
  wire [3:0] _GEN_194 = 7'h59 == _char_index_0_T_1[6:0] ? 4'h9 : _GEN_193; // @[CharOutput.scala 82:{21,21}]
  wire [3:0] _GEN_195 = 7'h5a == _char_index_0_T_1[6:0] ? 4'ha : _GEN_194; // @[CharOutput.scala 82:{21,21}]
  wire [3:0] _GEN_196 = 7'h5b == _char_index_0_T_1[6:0] ? 4'ha : _GEN_195; // @[CharOutput.scala 82:{21,21}]
  wire [3:0] _GEN_197 = 7'h5c == _char_index_0_T_1[6:0] ? 4'ha : _GEN_196; // @[CharOutput.scala 82:{21,21}]
  wire [3:0] _GEN_198 = 7'h5d == _char_index_0_T_1[6:0] ? 4'ha : _GEN_197; // @[CharOutput.scala 82:{21,21}]
  wire [3:0] _GEN_199 = 7'h5e == _char_index_0_T_1[6:0] ? 4'ha : _GEN_198; // @[CharOutput.scala 82:{21,21}]
  wire [3:0] _GEN_200 = 7'h5f == _char_index_0_T_1[6:0] ? 4'ha : _GEN_199; // @[CharOutput.scala 82:{21,21}]
  wire [3:0] _GEN_201 = 7'h60 == _char_index_0_T_1[6:0] ? 4'ha : _GEN_200; // @[CharOutput.scala 82:{21,21}]
  wire [3:0] _GEN_202 = 7'h61 == _char_index_0_T_1[6:0] ? 4'ha : _GEN_201; // @[CharOutput.scala 82:{21,21}]
  wire [3:0] _GEN_203 = 7'h62 == _char_index_0_T_1[6:0] ? 4'ha : _GEN_202; // @[CharOutput.scala 82:{21,21}]
  wire [3:0] _GEN_205 = 7'h1 == _char_index_0_T_1[6:0] ? 4'h1 : 4'h0; // @[CharOutput.scala 83:{19,19}]
  wire [3:0] _GEN_206 = 7'h2 == _char_index_0_T_1[6:0] ? 4'h2 : _GEN_205; // @[CharOutput.scala 83:{19,19}]
  wire [3:0] _GEN_207 = 7'h3 == _char_index_0_T_1[6:0] ? 4'h3 : _GEN_206; // @[CharOutput.scala 83:{19,19}]
  wire [3:0] _GEN_208 = 7'h4 == _char_index_0_T_1[6:0] ? 4'h4 : _GEN_207; // @[CharOutput.scala 83:{19,19}]
  wire [3:0] _GEN_209 = 7'h5 == _char_index_0_T_1[6:0] ? 4'h5 : _GEN_208; // @[CharOutput.scala 83:{19,19}]
  wire [3:0] _GEN_210 = 7'h6 == _char_index_0_T_1[6:0] ? 4'h6 : _GEN_209; // @[CharOutput.scala 83:{19,19}]
  wire [3:0] _GEN_211 = 7'h7 == _char_index_0_T_1[6:0] ? 4'h7 : _GEN_210; // @[CharOutput.scala 83:{19,19}]
  wire [3:0] _GEN_212 = 7'h8 == _char_index_0_T_1[6:0] ? 4'h8 : _GEN_211; // @[CharOutput.scala 83:{19,19}]
  wire [3:0] _GEN_213 = 7'h9 == _char_index_0_T_1[6:0] ? 4'h0 : _GEN_212; // @[CharOutput.scala 83:{19,19}]
  wire [3:0] _GEN_214 = 7'ha == _char_index_0_T_1[6:0] ? 4'h1 : _GEN_213; // @[CharOutput.scala 83:{19,19}]
  wire [3:0] _GEN_215 = 7'hb == _char_index_0_T_1[6:0] ? 4'h2 : _GEN_214; // @[CharOutput.scala 83:{19,19}]
  wire [3:0] _GEN_216 = 7'hc == _char_index_0_T_1[6:0] ? 4'h3 : _GEN_215; // @[CharOutput.scala 83:{19,19}]
  wire [3:0] _GEN_217 = 7'hd == _char_index_0_T_1[6:0] ? 4'h4 : _GEN_216; // @[CharOutput.scala 83:{19,19}]
  wire [3:0] _GEN_218 = 7'he == _char_index_0_T_1[6:0] ? 4'h5 : _GEN_217; // @[CharOutput.scala 83:{19,19}]
  wire [3:0] _GEN_219 = 7'hf == _char_index_0_T_1[6:0] ? 4'h6 : _GEN_218; // @[CharOutput.scala 83:{19,19}]
  wire [3:0] _GEN_220 = 7'h10 == _char_index_0_T_1[6:0] ? 4'h7 : _GEN_219; // @[CharOutput.scala 83:{19,19}]
  wire [3:0] _GEN_221 = 7'h11 == _char_index_0_T_1[6:0] ? 4'h8 : _GEN_220; // @[CharOutput.scala 83:{19,19}]
  wire [3:0] _GEN_222 = 7'h12 == _char_index_0_T_1[6:0] ? 4'h0 : _GEN_221; // @[CharOutput.scala 83:{19,19}]
  wire [3:0] _GEN_223 = 7'h13 == _char_index_0_T_1[6:0] ? 4'h1 : _GEN_222; // @[CharOutput.scala 83:{19,19}]
  wire [3:0] _GEN_224 = 7'h14 == _char_index_0_T_1[6:0] ? 4'h2 : _GEN_223; // @[CharOutput.scala 83:{19,19}]
  wire [3:0] _GEN_225 = 7'h15 == _char_index_0_T_1[6:0] ? 4'h3 : _GEN_224; // @[CharOutput.scala 83:{19,19}]
  wire [3:0] _GEN_226 = 7'h16 == _char_index_0_T_1[6:0] ? 4'h4 : _GEN_225; // @[CharOutput.scala 83:{19,19}]
  wire [3:0] _GEN_227 = 7'h17 == _char_index_0_T_1[6:0] ? 4'h5 : _GEN_226; // @[CharOutput.scala 83:{19,19}]
  wire [3:0] _GEN_228 = 7'h18 == _char_index_0_T_1[6:0] ? 4'h6 : _GEN_227; // @[CharOutput.scala 83:{19,19}]
  wire [3:0] _GEN_229 = 7'h19 == _char_index_0_T_1[6:0] ? 4'h7 : _GEN_228; // @[CharOutput.scala 83:{19,19}]
  wire [3:0] _GEN_230 = 7'h1a == _char_index_0_T_1[6:0] ? 4'h8 : _GEN_229; // @[CharOutput.scala 83:{19,19}]
  wire [3:0] _GEN_231 = 7'h1b == _char_index_0_T_1[6:0] ? 4'h0 : _GEN_230; // @[CharOutput.scala 83:{19,19}]
  wire [3:0] _GEN_232 = 7'h1c == _char_index_0_T_1[6:0] ? 4'h1 : _GEN_231; // @[CharOutput.scala 83:{19,19}]
  wire [3:0] _GEN_233 = 7'h1d == _char_index_0_T_1[6:0] ? 4'h2 : _GEN_232; // @[CharOutput.scala 83:{19,19}]
  wire [3:0] _GEN_234 = 7'h1e == _char_index_0_T_1[6:0] ? 4'h3 : _GEN_233; // @[CharOutput.scala 83:{19,19}]
  wire [3:0] _GEN_235 = 7'h1f == _char_index_0_T_1[6:0] ? 4'h4 : _GEN_234; // @[CharOutput.scala 83:{19,19}]
  wire [3:0] _GEN_236 = 7'h20 == _char_index_0_T_1[6:0] ? 4'h5 : _GEN_235; // @[CharOutput.scala 83:{19,19}]
  wire [3:0] _GEN_237 = 7'h21 == _char_index_0_T_1[6:0] ? 4'h6 : _GEN_236; // @[CharOutput.scala 83:{19,19}]
  wire [3:0] _GEN_238 = 7'h22 == _char_index_0_T_1[6:0] ? 4'h7 : _GEN_237; // @[CharOutput.scala 83:{19,19}]
  wire [3:0] _GEN_239 = 7'h23 == _char_index_0_T_1[6:0] ? 4'h8 : _GEN_238; // @[CharOutput.scala 83:{19,19}]
  wire [3:0] _GEN_240 = 7'h24 == _char_index_0_T_1[6:0] ? 4'h0 : _GEN_239; // @[CharOutput.scala 83:{19,19}]
  wire [3:0] _GEN_241 = 7'h25 == _char_index_0_T_1[6:0] ? 4'h1 : _GEN_240; // @[CharOutput.scala 83:{19,19}]
  wire [3:0] _GEN_242 = 7'h26 == _char_index_0_T_1[6:0] ? 4'h2 : _GEN_241; // @[CharOutput.scala 83:{19,19}]
  wire [3:0] _GEN_243 = 7'h27 == _char_index_0_T_1[6:0] ? 4'h3 : _GEN_242; // @[CharOutput.scala 83:{19,19}]
  wire [3:0] _GEN_244 = 7'h28 == _char_index_0_T_1[6:0] ? 4'h4 : _GEN_243; // @[CharOutput.scala 83:{19,19}]
  wire [3:0] _GEN_245 = 7'h29 == _char_index_0_T_1[6:0] ? 4'h5 : _GEN_244; // @[CharOutput.scala 83:{19,19}]
  wire [3:0] _GEN_246 = 7'h2a == _char_index_0_T_1[6:0] ? 4'h6 : _GEN_245; // @[CharOutput.scala 83:{19,19}]
  wire [3:0] _GEN_247 = 7'h2b == _char_index_0_T_1[6:0] ? 4'h7 : _GEN_246; // @[CharOutput.scala 83:{19,19}]
  wire [3:0] _GEN_248 = 7'h2c == _char_index_0_T_1[6:0] ? 4'h8 : _GEN_247; // @[CharOutput.scala 83:{19,19}]
  wire [3:0] _GEN_249 = 7'h2d == _char_index_0_T_1[6:0] ? 4'h0 : _GEN_248; // @[CharOutput.scala 83:{19,19}]
  wire [3:0] _GEN_250 = 7'h2e == _char_index_0_T_1[6:0] ? 4'h1 : _GEN_249; // @[CharOutput.scala 83:{19,19}]
  wire [3:0] _GEN_251 = 7'h2f == _char_index_0_T_1[6:0] ? 4'h2 : _GEN_250; // @[CharOutput.scala 83:{19,19}]
  wire [3:0] _GEN_252 = 7'h30 == _char_index_0_T_1[6:0] ? 4'h3 : _GEN_251; // @[CharOutput.scala 83:{19,19}]
  wire [3:0] _GEN_253 = 7'h31 == _char_index_0_T_1[6:0] ? 4'h4 : _GEN_252; // @[CharOutput.scala 83:{19,19}]
  wire [3:0] _GEN_254 = 7'h32 == _char_index_0_T_1[6:0] ? 4'h5 : _GEN_253; // @[CharOutput.scala 83:{19,19}]
  wire [3:0] _GEN_255 = 7'h33 == _char_index_0_T_1[6:0] ? 4'h6 : _GEN_254; // @[CharOutput.scala 83:{19,19}]
  wire [3:0] _GEN_256 = 7'h34 == _char_index_0_T_1[6:0] ? 4'h7 : _GEN_255; // @[CharOutput.scala 83:{19,19}]
  wire [3:0] _GEN_257 = 7'h35 == _char_index_0_T_1[6:0] ? 4'h8 : _GEN_256; // @[CharOutput.scala 83:{19,19}]
  wire [3:0] _GEN_258 = 7'h36 == _char_index_0_T_1[6:0] ? 4'h0 : _GEN_257; // @[CharOutput.scala 83:{19,19}]
  wire [3:0] _GEN_259 = 7'h37 == _char_index_0_T_1[6:0] ? 4'h1 : _GEN_258; // @[CharOutput.scala 83:{19,19}]
  wire [3:0] _GEN_260 = 7'h38 == _char_index_0_T_1[6:0] ? 4'h2 : _GEN_259; // @[CharOutput.scala 83:{19,19}]
  wire [3:0] _GEN_261 = 7'h39 == _char_index_0_T_1[6:0] ? 4'h3 : _GEN_260; // @[CharOutput.scala 83:{19,19}]
  wire [3:0] _GEN_262 = 7'h3a == _char_index_0_T_1[6:0] ? 4'h4 : _GEN_261; // @[CharOutput.scala 83:{19,19}]
  wire [3:0] _GEN_263 = 7'h3b == _char_index_0_T_1[6:0] ? 4'h5 : _GEN_262; // @[CharOutput.scala 83:{19,19}]
  wire [3:0] _GEN_264 = 7'h3c == _char_index_0_T_1[6:0] ? 4'h6 : _GEN_263; // @[CharOutput.scala 83:{19,19}]
  wire [3:0] _GEN_265 = 7'h3d == _char_index_0_T_1[6:0] ? 4'h7 : _GEN_264; // @[CharOutput.scala 83:{19,19}]
  wire [3:0] _GEN_266 = 7'h3e == _char_index_0_T_1[6:0] ? 4'h8 : _GEN_265; // @[CharOutput.scala 83:{19,19}]
  wire [3:0] _GEN_267 = 7'h3f == _char_index_0_T_1[6:0] ? 4'h0 : _GEN_266; // @[CharOutput.scala 83:{19,19}]
  wire [3:0] _GEN_268 = 7'h40 == _char_index_0_T_1[6:0] ? 4'h1 : _GEN_267; // @[CharOutput.scala 83:{19,19}]
  wire [3:0] _GEN_269 = 7'h41 == _char_index_0_T_1[6:0] ? 4'h2 : _GEN_268; // @[CharOutput.scala 83:{19,19}]
  wire [3:0] _GEN_270 = 7'h42 == _char_index_0_T_1[6:0] ? 4'h3 : _GEN_269; // @[CharOutput.scala 83:{19,19}]
  wire [3:0] _GEN_271 = 7'h43 == _char_index_0_T_1[6:0] ? 4'h4 : _GEN_270; // @[CharOutput.scala 83:{19,19}]
  wire [3:0] _GEN_272 = 7'h44 == _char_index_0_T_1[6:0] ? 4'h5 : _GEN_271; // @[CharOutput.scala 83:{19,19}]
  wire [3:0] _GEN_273 = 7'h45 == _char_index_0_T_1[6:0] ? 4'h6 : _GEN_272; // @[CharOutput.scala 83:{19,19}]
  wire [3:0] _GEN_274 = 7'h46 == _char_index_0_T_1[6:0] ? 4'h7 : _GEN_273; // @[CharOutput.scala 83:{19,19}]
  wire [3:0] _GEN_275 = 7'h47 == _char_index_0_T_1[6:0] ? 4'h8 : _GEN_274; // @[CharOutput.scala 83:{19,19}]
  wire [3:0] _GEN_276 = 7'h48 == _char_index_0_T_1[6:0] ? 4'h0 : _GEN_275; // @[CharOutput.scala 83:{19,19}]
  wire [3:0] _GEN_277 = 7'h49 == _char_index_0_T_1[6:0] ? 4'h1 : _GEN_276; // @[CharOutput.scala 83:{19,19}]
  wire [3:0] _GEN_278 = 7'h4a == _char_index_0_T_1[6:0] ? 4'h2 : _GEN_277; // @[CharOutput.scala 83:{19,19}]
  wire [3:0] _GEN_279 = 7'h4b == _char_index_0_T_1[6:0] ? 4'h3 : _GEN_278; // @[CharOutput.scala 83:{19,19}]
  wire [3:0] _GEN_280 = 7'h4c == _char_index_0_T_1[6:0] ? 4'h4 : _GEN_279; // @[CharOutput.scala 83:{19,19}]
  wire [3:0] _GEN_281 = 7'h4d == _char_index_0_T_1[6:0] ? 4'h5 : _GEN_280; // @[CharOutput.scala 83:{19,19}]
  wire [3:0] _GEN_282 = 7'h4e == _char_index_0_T_1[6:0] ? 4'h6 : _GEN_281; // @[CharOutput.scala 83:{19,19}]
  wire [3:0] _GEN_283 = 7'h4f == _char_index_0_T_1[6:0] ? 4'h7 : _GEN_282; // @[CharOutput.scala 83:{19,19}]
  wire [3:0] _GEN_284 = 7'h50 == _char_index_0_T_1[6:0] ? 4'h8 : _GEN_283; // @[CharOutput.scala 83:{19,19}]
  wire [3:0] _GEN_285 = 7'h51 == _char_index_0_T_1[6:0] ? 4'h0 : _GEN_284; // @[CharOutput.scala 83:{19,19}]
  wire [3:0] _GEN_286 = 7'h52 == _char_index_0_T_1[6:0] ? 4'h1 : _GEN_285; // @[CharOutput.scala 83:{19,19}]
  wire [3:0] _GEN_287 = 7'h53 == _char_index_0_T_1[6:0] ? 4'h2 : _GEN_286; // @[CharOutput.scala 83:{19,19}]
  wire [3:0] _GEN_288 = 7'h54 == _char_index_0_T_1[6:0] ? 4'h3 : _GEN_287; // @[CharOutput.scala 83:{19,19}]
  wire [3:0] _GEN_289 = 7'h55 == _char_index_0_T_1[6:0] ? 4'h4 : _GEN_288; // @[CharOutput.scala 83:{19,19}]
  wire [3:0] _GEN_290 = 7'h56 == _char_index_0_T_1[6:0] ? 4'h5 : _GEN_289; // @[CharOutput.scala 83:{19,19}]
  wire [3:0] _GEN_291 = 7'h57 == _char_index_0_T_1[6:0] ? 4'h6 : _GEN_290; // @[CharOutput.scala 83:{19,19}]
  wire [3:0] _GEN_292 = 7'h58 == _char_index_0_T_1[6:0] ? 4'h7 : _GEN_291; // @[CharOutput.scala 83:{19,19}]
  wire [3:0] _GEN_293 = 7'h59 == _char_index_0_T_1[6:0] ? 4'h8 : _GEN_292; // @[CharOutput.scala 83:{19,19}]
  wire [3:0] _GEN_294 = 7'h5a == _char_index_0_T_1[6:0] ? 4'h0 : _GEN_293; // @[CharOutput.scala 83:{19,19}]
  wire [3:0] _GEN_295 = 7'h5b == _char_index_0_T_1[6:0] ? 4'h1 : _GEN_294; // @[CharOutput.scala 83:{19,19}]
  wire [3:0] _GEN_296 = 7'h5c == _char_index_0_T_1[6:0] ? 4'h2 : _GEN_295; // @[CharOutput.scala 83:{19,19}]
  wire [3:0] _GEN_297 = 7'h5d == _char_index_0_T_1[6:0] ? 4'h3 : _GEN_296; // @[CharOutput.scala 83:{19,19}]
  wire [3:0] _GEN_298 = 7'h5e == _char_index_0_T_1[6:0] ? 4'h4 : _GEN_297; // @[CharOutput.scala 83:{19,19}]
  wire [3:0] _GEN_299 = 7'h5f == _char_index_0_T_1[6:0] ? 4'h5 : _GEN_298; // @[CharOutput.scala 83:{19,19}]
  wire [3:0] _GEN_300 = 7'h60 == _char_index_0_T_1[6:0] ? 4'h6 : _GEN_299; // @[CharOutput.scala 83:{19,19}]
  wire [3:0] _GEN_301 = 7'h61 == _char_index_0_T_1[6:0] ? 4'h7 : _GEN_300; // @[CharOutput.scala 83:{19,19}]
  wire [3:0] _GEN_302 = 7'h62 == _char_index_0_T_1[6:0] ? 4'h8 : _GEN_301; // @[CharOutput.scala 83:{19,19}]
  wire [3:0] char_index_0 = in_area_h_0 ? _GEN_203 : 4'h0; // @[CharOutput.scala 81:23 82:21 85:21]
  wire [3:0] char_col_0 = in_area_h_0 ? _GEN_302 : 4'h0; // @[CharOutput.scala 81:23 83:19 86:19]
  wire [10:0] _char_row_0_T_1 = io_v_cnt - char_area_ytop_0; // @[CharOutput.scala 89:31]
  wire [10:0] _GEN_305 = in_area_v_0 ? _char_row_0_T_1 : 11'h0; // @[CharOutput.scala 88:23 89:19 91:19]
  wire [10:0] _char_index_1_T_1 = io_h_cnt - io_rect_xleft_1; // @[CharOutput.scala 82:48]
  wire [3:0] _GEN_315 = 7'h9 == _char_index_1_T_1[6:0] ? 4'h1 : 4'h0; // @[CharOutput.scala 82:{21,21}]
  wire [3:0] _GEN_316 = 7'ha == _char_index_1_T_1[6:0] ? 4'h1 : _GEN_315; // @[CharOutput.scala 82:{21,21}]
  wire [3:0] _GEN_317 = 7'hb == _char_index_1_T_1[6:0] ? 4'h1 : _GEN_316; // @[CharOutput.scala 82:{21,21}]
  wire [3:0] _GEN_318 = 7'hc == _char_index_1_T_1[6:0] ? 4'h1 : _GEN_317; // @[CharOutput.scala 82:{21,21}]
  wire [3:0] _GEN_319 = 7'hd == _char_index_1_T_1[6:0] ? 4'h1 : _GEN_318; // @[CharOutput.scala 82:{21,21}]
  wire [3:0] _GEN_320 = 7'he == _char_index_1_T_1[6:0] ? 4'h1 : _GEN_319; // @[CharOutput.scala 82:{21,21}]
  wire [3:0] _GEN_321 = 7'hf == _char_index_1_T_1[6:0] ? 4'h1 : _GEN_320; // @[CharOutput.scala 82:{21,21}]
  wire [3:0] _GEN_322 = 7'h10 == _char_index_1_T_1[6:0] ? 4'h1 : _GEN_321; // @[CharOutput.scala 82:{21,21}]
  wire [3:0] _GEN_323 = 7'h11 == _char_index_1_T_1[6:0] ? 4'h1 : _GEN_322; // @[CharOutput.scala 82:{21,21}]
  wire [3:0] _GEN_324 = 7'h12 == _char_index_1_T_1[6:0] ? 4'h2 : _GEN_323; // @[CharOutput.scala 82:{21,21}]
  wire [3:0] _GEN_325 = 7'h13 == _char_index_1_T_1[6:0] ? 4'h2 : _GEN_324; // @[CharOutput.scala 82:{21,21}]
  wire [3:0] _GEN_326 = 7'h14 == _char_index_1_T_1[6:0] ? 4'h2 : _GEN_325; // @[CharOutput.scala 82:{21,21}]
  wire [3:0] _GEN_327 = 7'h15 == _char_index_1_T_1[6:0] ? 4'h2 : _GEN_326; // @[CharOutput.scala 82:{21,21}]
  wire [3:0] _GEN_328 = 7'h16 == _char_index_1_T_1[6:0] ? 4'h2 : _GEN_327; // @[CharOutput.scala 82:{21,21}]
  wire [3:0] _GEN_329 = 7'h17 == _char_index_1_T_1[6:0] ? 4'h2 : _GEN_328; // @[CharOutput.scala 82:{21,21}]
  wire [3:0] _GEN_330 = 7'h18 == _char_index_1_T_1[6:0] ? 4'h2 : _GEN_329; // @[CharOutput.scala 82:{21,21}]
  wire [3:0] _GEN_331 = 7'h19 == _char_index_1_T_1[6:0] ? 4'h2 : _GEN_330; // @[CharOutput.scala 82:{21,21}]
  wire [3:0] _GEN_332 = 7'h1a == _char_index_1_T_1[6:0] ? 4'h2 : _GEN_331; // @[CharOutput.scala 82:{21,21}]
  wire [3:0] _GEN_333 = 7'h1b == _char_index_1_T_1[6:0] ? 4'h3 : _GEN_332; // @[CharOutput.scala 82:{21,21}]
  wire [3:0] _GEN_334 = 7'h1c == _char_index_1_T_1[6:0] ? 4'h3 : _GEN_333; // @[CharOutput.scala 82:{21,21}]
  wire [3:0] _GEN_335 = 7'h1d == _char_index_1_T_1[6:0] ? 4'h3 : _GEN_334; // @[CharOutput.scala 82:{21,21}]
  wire [3:0] _GEN_336 = 7'h1e == _char_index_1_T_1[6:0] ? 4'h3 : _GEN_335; // @[CharOutput.scala 82:{21,21}]
  wire [3:0] _GEN_337 = 7'h1f == _char_index_1_T_1[6:0] ? 4'h3 : _GEN_336; // @[CharOutput.scala 82:{21,21}]
  wire [3:0] _GEN_338 = 7'h20 == _char_index_1_T_1[6:0] ? 4'h3 : _GEN_337; // @[CharOutput.scala 82:{21,21}]
  wire [3:0] _GEN_339 = 7'h21 == _char_index_1_T_1[6:0] ? 4'h3 : _GEN_338; // @[CharOutput.scala 82:{21,21}]
  wire [3:0] _GEN_340 = 7'h22 == _char_index_1_T_1[6:0] ? 4'h3 : _GEN_339; // @[CharOutput.scala 82:{21,21}]
  wire [3:0] _GEN_341 = 7'h23 == _char_index_1_T_1[6:0] ? 4'h3 : _GEN_340; // @[CharOutput.scala 82:{21,21}]
  wire [3:0] _GEN_342 = 7'h24 == _char_index_1_T_1[6:0] ? 4'h4 : _GEN_341; // @[CharOutput.scala 82:{21,21}]
  wire [3:0] _GEN_343 = 7'h25 == _char_index_1_T_1[6:0] ? 4'h4 : _GEN_342; // @[CharOutput.scala 82:{21,21}]
  wire [3:0] _GEN_344 = 7'h26 == _char_index_1_T_1[6:0] ? 4'h4 : _GEN_343; // @[CharOutput.scala 82:{21,21}]
  wire [3:0] _GEN_345 = 7'h27 == _char_index_1_T_1[6:0] ? 4'h4 : _GEN_344; // @[CharOutput.scala 82:{21,21}]
  wire [3:0] _GEN_346 = 7'h28 == _char_index_1_T_1[6:0] ? 4'h4 : _GEN_345; // @[CharOutput.scala 82:{21,21}]
  wire [3:0] _GEN_347 = 7'h29 == _char_index_1_T_1[6:0] ? 4'h4 : _GEN_346; // @[CharOutput.scala 82:{21,21}]
  wire [3:0] _GEN_348 = 7'h2a == _char_index_1_T_1[6:0] ? 4'h4 : _GEN_347; // @[CharOutput.scala 82:{21,21}]
  wire [3:0] _GEN_349 = 7'h2b == _char_index_1_T_1[6:0] ? 4'h4 : _GEN_348; // @[CharOutput.scala 82:{21,21}]
  wire [3:0] _GEN_350 = 7'h2c == _char_index_1_T_1[6:0] ? 4'h4 : _GEN_349; // @[CharOutput.scala 82:{21,21}]
  wire [3:0] _GEN_351 = 7'h2d == _char_index_1_T_1[6:0] ? 4'h5 : _GEN_350; // @[CharOutput.scala 82:{21,21}]
  wire [3:0] _GEN_352 = 7'h2e == _char_index_1_T_1[6:0] ? 4'h5 : _GEN_351; // @[CharOutput.scala 82:{21,21}]
  wire [3:0] _GEN_353 = 7'h2f == _char_index_1_T_1[6:0] ? 4'h5 : _GEN_352; // @[CharOutput.scala 82:{21,21}]
  wire [3:0] _GEN_354 = 7'h30 == _char_index_1_T_1[6:0] ? 4'h5 : _GEN_353; // @[CharOutput.scala 82:{21,21}]
  wire [3:0] _GEN_355 = 7'h31 == _char_index_1_T_1[6:0] ? 4'h5 : _GEN_354; // @[CharOutput.scala 82:{21,21}]
  wire [3:0] _GEN_356 = 7'h32 == _char_index_1_T_1[6:0] ? 4'h5 : _GEN_355; // @[CharOutput.scala 82:{21,21}]
  wire [3:0] _GEN_357 = 7'h33 == _char_index_1_T_1[6:0] ? 4'h5 : _GEN_356; // @[CharOutput.scala 82:{21,21}]
  wire [3:0] _GEN_358 = 7'h34 == _char_index_1_T_1[6:0] ? 4'h5 : _GEN_357; // @[CharOutput.scala 82:{21,21}]
  wire [3:0] _GEN_359 = 7'h35 == _char_index_1_T_1[6:0] ? 4'h5 : _GEN_358; // @[CharOutput.scala 82:{21,21}]
  wire [3:0] _GEN_360 = 7'h36 == _char_index_1_T_1[6:0] ? 4'h6 : _GEN_359; // @[CharOutput.scala 82:{21,21}]
  wire [3:0] _GEN_361 = 7'h37 == _char_index_1_T_1[6:0] ? 4'h6 : _GEN_360; // @[CharOutput.scala 82:{21,21}]
  wire [3:0] _GEN_362 = 7'h38 == _char_index_1_T_1[6:0] ? 4'h6 : _GEN_361; // @[CharOutput.scala 82:{21,21}]
  wire [3:0] _GEN_363 = 7'h39 == _char_index_1_T_1[6:0] ? 4'h6 : _GEN_362; // @[CharOutput.scala 82:{21,21}]
  wire [3:0] _GEN_364 = 7'h3a == _char_index_1_T_1[6:0] ? 4'h6 : _GEN_363; // @[CharOutput.scala 82:{21,21}]
  wire [3:0] _GEN_365 = 7'h3b == _char_index_1_T_1[6:0] ? 4'h6 : _GEN_364; // @[CharOutput.scala 82:{21,21}]
  wire [3:0] _GEN_366 = 7'h3c == _char_index_1_T_1[6:0] ? 4'h6 : _GEN_365; // @[CharOutput.scala 82:{21,21}]
  wire [3:0] _GEN_367 = 7'h3d == _char_index_1_T_1[6:0] ? 4'h6 : _GEN_366; // @[CharOutput.scala 82:{21,21}]
  wire [3:0] _GEN_368 = 7'h3e == _char_index_1_T_1[6:0] ? 4'h6 : _GEN_367; // @[CharOutput.scala 82:{21,21}]
  wire [3:0] _GEN_369 = 7'h3f == _char_index_1_T_1[6:0] ? 4'h7 : _GEN_368; // @[CharOutput.scala 82:{21,21}]
  wire [3:0] _GEN_370 = 7'h40 == _char_index_1_T_1[6:0] ? 4'h7 : _GEN_369; // @[CharOutput.scala 82:{21,21}]
  wire [3:0] _GEN_371 = 7'h41 == _char_index_1_T_1[6:0] ? 4'h7 : _GEN_370; // @[CharOutput.scala 82:{21,21}]
  wire [3:0] _GEN_372 = 7'h42 == _char_index_1_T_1[6:0] ? 4'h7 : _GEN_371; // @[CharOutput.scala 82:{21,21}]
  wire [3:0] _GEN_373 = 7'h43 == _char_index_1_T_1[6:0] ? 4'h7 : _GEN_372; // @[CharOutput.scala 82:{21,21}]
  wire [3:0] _GEN_374 = 7'h44 == _char_index_1_T_1[6:0] ? 4'h7 : _GEN_373; // @[CharOutput.scala 82:{21,21}]
  wire [3:0] _GEN_375 = 7'h45 == _char_index_1_T_1[6:0] ? 4'h7 : _GEN_374; // @[CharOutput.scala 82:{21,21}]
  wire [3:0] _GEN_376 = 7'h46 == _char_index_1_T_1[6:0] ? 4'h7 : _GEN_375; // @[CharOutput.scala 82:{21,21}]
  wire [3:0] _GEN_377 = 7'h47 == _char_index_1_T_1[6:0] ? 4'h7 : _GEN_376; // @[CharOutput.scala 82:{21,21}]
  wire [3:0] _GEN_378 = 7'h48 == _char_index_1_T_1[6:0] ? 4'h8 : _GEN_377; // @[CharOutput.scala 82:{21,21}]
  wire [3:0] _GEN_379 = 7'h49 == _char_index_1_T_1[6:0] ? 4'h8 : _GEN_378; // @[CharOutput.scala 82:{21,21}]
  wire [3:0] _GEN_380 = 7'h4a == _char_index_1_T_1[6:0] ? 4'h8 : _GEN_379; // @[CharOutput.scala 82:{21,21}]
  wire [3:0] _GEN_381 = 7'h4b == _char_index_1_T_1[6:0] ? 4'h8 : _GEN_380; // @[CharOutput.scala 82:{21,21}]
  wire [3:0] _GEN_382 = 7'h4c == _char_index_1_T_1[6:0] ? 4'h8 : _GEN_381; // @[CharOutput.scala 82:{21,21}]
  wire [3:0] _GEN_383 = 7'h4d == _char_index_1_T_1[6:0] ? 4'h8 : _GEN_382; // @[CharOutput.scala 82:{21,21}]
  wire [3:0] _GEN_384 = 7'h4e == _char_index_1_T_1[6:0] ? 4'h8 : _GEN_383; // @[CharOutput.scala 82:{21,21}]
  wire [3:0] _GEN_385 = 7'h4f == _char_index_1_T_1[6:0] ? 4'h8 : _GEN_384; // @[CharOutput.scala 82:{21,21}]
  wire [3:0] _GEN_386 = 7'h50 == _char_index_1_T_1[6:0] ? 4'h8 : _GEN_385; // @[CharOutput.scala 82:{21,21}]
  wire [3:0] _GEN_387 = 7'h51 == _char_index_1_T_1[6:0] ? 4'h9 : _GEN_386; // @[CharOutput.scala 82:{21,21}]
  wire [3:0] _GEN_388 = 7'h52 == _char_index_1_T_1[6:0] ? 4'h9 : _GEN_387; // @[CharOutput.scala 82:{21,21}]
  wire [3:0] _GEN_389 = 7'h53 == _char_index_1_T_1[6:0] ? 4'h9 : _GEN_388; // @[CharOutput.scala 82:{21,21}]
  wire [3:0] _GEN_390 = 7'h54 == _char_index_1_T_1[6:0] ? 4'h9 : _GEN_389; // @[CharOutput.scala 82:{21,21}]
  wire [3:0] _GEN_391 = 7'h55 == _char_index_1_T_1[6:0] ? 4'h9 : _GEN_390; // @[CharOutput.scala 82:{21,21}]
  wire [3:0] _GEN_392 = 7'h56 == _char_index_1_T_1[6:0] ? 4'h9 : _GEN_391; // @[CharOutput.scala 82:{21,21}]
  wire [3:0] _GEN_393 = 7'h57 == _char_index_1_T_1[6:0] ? 4'h9 : _GEN_392; // @[CharOutput.scala 82:{21,21}]
  wire [3:0] _GEN_394 = 7'h58 == _char_index_1_T_1[6:0] ? 4'h9 : _GEN_393; // @[CharOutput.scala 82:{21,21}]
  wire [3:0] _GEN_395 = 7'h59 == _char_index_1_T_1[6:0] ? 4'h9 : _GEN_394; // @[CharOutput.scala 82:{21,21}]
  wire [3:0] _GEN_396 = 7'h5a == _char_index_1_T_1[6:0] ? 4'ha : _GEN_395; // @[CharOutput.scala 82:{21,21}]
  wire [3:0] _GEN_397 = 7'h5b == _char_index_1_T_1[6:0] ? 4'ha : _GEN_396; // @[CharOutput.scala 82:{21,21}]
  wire [3:0] _GEN_398 = 7'h5c == _char_index_1_T_1[6:0] ? 4'ha : _GEN_397; // @[CharOutput.scala 82:{21,21}]
  wire [3:0] _GEN_399 = 7'h5d == _char_index_1_T_1[6:0] ? 4'ha : _GEN_398; // @[CharOutput.scala 82:{21,21}]
  wire [3:0] _GEN_400 = 7'h5e == _char_index_1_T_1[6:0] ? 4'ha : _GEN_399; // @[CharOutput.scala 82:{21,21}]
  wire [3:0] _GEN_401 = 7'h5f == _char_index_1_T_1[6:0] ? 4'ha : _GEN_400; // @[CharOutput.scala 82:{21,21}]
  wire [3:0] _GEN_402 = 7'h60 == _char_index_1_T_1[6:0] ? 4'ha : _GEN_401; // @[CharOutput.scala 82:{21,21}]
  wire [3:0] _GEN_403 = 7'h61 == _char_index_1_T_1[6:0] ? 4'ha : _GEN_402; // @[CharOutput.scala 82:{21,21}]
  wire [3:0] _GEN_404 = 7'h62 == _char_index_1_T_1[6:0] ? 4'ha : _GEN_403; // @[CharOutput.scala 82:{21,21}]
  wire [3:0] _GEN_406 = 7'h1 == _char_index_1_T_1[6:0] ? 4'h1 : 4'h0; // @[CharOutput.scala 83:{19,19}]
  wire [3:0] _GEN_407 = 7'h2 == _char_index_1_T_1[6:0] ? 4'h2 : _GEN_406; // @[CharOutput.scala 83:{19,19}]
  wire [3:0] _GEN_408 = 7'h3 == _char_index_1_T_1[6:0] ? 4'h3 : _GEN_407; // @[CharOutput.scala 83:{19,19}]
  wire [3:0] _GEN_409 = 7'h4 == _char_index_1_T_1[6:0] ? 4'h4 : _GEN_408; // @[CharOutput.scala 83:{19,19}]
  wire [3:0] _GEN_410 = 7'h5 == _char_index_1_T_1[6:0] ? 4'h5 : _GEN_409; // @[CharOutput.scala 83:{19,19}]
  wire [3:0] _GEN_411 = 7'h6 == _char_index_1_T_1[6:0] ? 4'h6 : _GEN_410; // @[CharOutput.scala 83:{19,19}]
  wire [3:0] _GEN_412 = 7'h7 == _char_index_1_T_1[6:0] ? 4'h7 : _GEN_411; // @[CharOutput.scala 83:{19,19}]
  wire [3:0] _GEN_413 = 7'h8 == _char_index_1_T_1[6:0] ? 4'h8 : _GEN_412; // @[CharOutput.scala 83:{19,19}]
  wire [3:0] _GEN_414 = 7'h9 == _char_index_1_T_1[6:0] ? 4'h0 : _GEN_413; // @[CharOutput.scala 83:{19,19}]
  wire [3:0] _GEN_415 = 7'ha == _char_index_1_T_1[6:0] ? 4'h1 : _GEN_414; // @[CharOutput.scala 83:{19,19}]
  wire [3:0] _GEN_416 = 7'hb == _char_index_1_T_1[6:0] ? 4'h2 : _GEN_415; // @[CharOutput.scala 83:{19,19}]
  wire [3:0] _GEN_417 = 7'hc == _char_index_1_T_1[6:0] ? 4'h3 : _GEN_416; // @[CharOutput.scala 83:{19,19}]
  wire [3:0] _GEN_418 = 7'hd == _char_index_1_T_1[6:0] ? 4'h4 : _GEN_417; // @[CharOutput.scala 83:{19,19}]
  wire [3:0] _GEN_419 = 7'he == _char_index_1_T_1[6:0] ? 4'h5 : _GEN_418; // @[CharOutput.scala 83:{19,19}]
  wire [3:0] _GEN_420 = 7'hf == _char_index_1_T_1[6:0] ? 4'h6 : _GEN_419; // @[CharOutput.scala 83:{19,19}]
  wire [3:0] _GEN_421 = 7'h10 == _char_index_1_T_1[6:0] ? 4'h7 : _GEN_420; // @[CharOutput.scala 83:{19,19}]
  wire [3:0] _GEN_422 = 7'h11 == _char_index_1_T_1[6:0] ? 4'h8 : _GEN_421; // @[CharOutput.scala 83:{19,19}]
  wire [3:0] _GEN_423 = 7'h12 == _char_index_1_T_1[6:0] ? 4'h0 : _GEN_422; // @[CharOutput.scala 83:{19,19}]
  wire [3:0] _GEN_424 = 7'h13 == _char_index_1_T_1[6:0] ? 4'h1 : _GEN_423; // @[CharOutput.scala 83:{19,19}]
  wire [3:0] _GEN_425 = 7'h14 == _char_index_1_T_1[6:0] ? 4'h2 : _GEN_424; // @[CharOutput.scala 83:{19,19}]
  wire [3:0] _GEN_426 = 7'h15 == _char_index_1_T_1[6:0] ? 4'h3 : _GEN_425; // @[CharOutput.scala 83:{19,19}]
  wire [3:0] _GEN_427 = 7'h16 == _char_index_1_T_1[6:0] ? 4'h4 : _GEN_426; // @[CharOutput.scala 83:{19,19}]
  wire [3:0] _GEN_428 = 7'h17 == _char_index_1_T_1[6:0] ? 4'h5 : _GEN_427; // @[CharOutput.scala 83:{19,19}]
  wire [3:0] _GEN_429 = 7'h18 == _char_index_1_T_1[6:0] ? 4'h6 : _GEN_428; // @[CharOutput.scala 83:{19,19}]
  wire [3:0] _GEN_430 = 7'h19 == _char_index_1_T_1[6:0] ? 4'h7 : _GEN_429; // @[CharOutput.scala 83:{19,19}]
  wire [3:0] _GEN_431 = 7'h1a == _char_index_1_T_1[6:0] ? 4'h8 : _GEN_430; // @[CharOutput.scala 83:{19,19}]
  wire [3:0] _GEN_432 = 7'h1b == _char_index_1_T_1[6:0] ? 4'h0 : _GEN_431; // @[CharOutput.scala 83:{19,19}]
  wire [3:0] _GEN_433 = 7'h1c == _char_index_1_T_1[6:0] ? 4'h1 : _GEN_432; // @[CharOutput.scala 83:{19,19}]
  wire [3:0] _GEN_434 = 7'h1d == _char_index_1_T_1[6:0] ? 4'h2 : _GEN_433; // @[CharOutput.scala 83:{19,19}]
  wire [3:0] _GEN_435 = 7'h1e == _char_index_1_T_1[6:0] ? 4'h3 : _GEN_434; // @[CharOutput.scala 83:{19,19}]
  wire [3:0] _GEN_436 = 7'h1f == _char_index_1_T_1[6:0] ? 4'h4 : _GEN_435; // @[CharOutput.scala 83:{19,19}]
  wire [3:0] _GEN_437 = 7'h20 == _char_index_1_T_1[6:0] ? 4'h5 : _GEN_436; // @[CharOutput.scala 83:{19,19}]
  wire [3:0] _GEN_438 = 7'h21 == _char_index_1_T_1[6:0] ? 4'h6 : _GEN_437; // @[CharOutput.scala 83:{19,19}]
  wire [3:0] _GEN_439 = 7'h22 == _char_index_1_T_1[6:0] ? 4'h7 : _GEN_438; // @[CharOutput.scala 83:{19,19}]
  wire [3:0] _GEN_440 = 7'h23 == _char_index_1_T_1[6:0] ? 4'h8 : _GEN_439; // @[CharOutput.scala 83:{19,19}]
  wire [3:0] _GEN_441 = 7'h24 == _char_index_1_T_1[6:0] ? 4'h0 : _GEN_440; // @[CharOutput.scala 83:{19,19}]
  wire [3:0] _GEN_442 = 7'h25 == _char_index_1_T_1[6:0] ? 4'h1 : _GEN_441; // @[CharOutput.scala 83:{19,19}]
  wire [3:0] _GEN_443 = 7'h26 == _char_index_1_T_1[6:0] ? 4'h2 : _GEN_442; // @[CharOutput.scala 83:{19,19}]
  wire [3:0] _GEN_444 = 7'h27 == _char_index_1_T_1[6:0] ? 4'h3 : _GEN_443; // @[CharOutput.scala 83:{19,19}]
  wire [3:0] _GEN_445 = 7'h28 == _char_index_1_T_1[6:0] ? 4'h4 : _GEN_444; // @[CharOutput.scala 83:{19,19}]
  wire [3:0] _GEN_446 = 7'h29 == _char_index_1_T_1[6:0] ? 4'h5 : _GEN_445; // @[CharOutput.scala 83:{19,19}]
  wire [3:0] _GEN_447 = 7'h2a == _char_index_1_T_1[6:0] ? 4'h6 : _GEN_446; // @[CharOutput.scala 83:{19,19}]
  wire [3:0] _GEN_448 = 7'h2b == _char_index_1_T_1[6:0] ? 4'h7 : _GEN_447; // @[CharOutput.scala 83:{19,19}]
  wire [3:0] _GEN_449 = 7'h2c == _char_index_1_T_1[6:0] ? 4'h8 : _GEN_448; // @[CharOutput.scala 83:{19,19}]
  wire [3:0] _GEN_450 = 7'h2d == _char_index_1_T_1[6:0] ? 4'h0 : _GEN_449; // @[CharOutput.scala 83:{19,19}]
  wire [3:0] _GEN_451 = 7'h2e == _char_index_1_T_1[6:0] ? 4'h1 : _GEN_450; // @[CharOutput.scala 83:{19,19}]
  wire [3:0] _GEN_452 = 7'h2f == _char_index_1_T_1[6:0] ? 4'h2 : _GEN_451; // @[CharOutput.scala 83:{19,19}]
  wire [3:0] _GEN_453 = 7'h30 == _char_index_1_T_1[6:0] ? 4'h3 : _GEN_452; // @[CharOutput.scala 83:{19,19}]
  wire [3:0] _GEN_454 = 7'h31 == _char_index_1_T_1[6:0] ? 4'h4 : _GEN_453; // @[CharOutput.scala 83:{19,19}]
  wire [3:0] _GEN_455 = 7'h32 == _char_index_1_T_1[6:0] ? 4'h5 : _GEN_454; // @[CharOutput.scala 83:{19,19}]
  wire [3:0] _GEN_456 = 7'h33 == _char_index_1_T_1[6:0] ? 4'h6 : _GEN_455; // @[CharOutput.scala 83:{19,19}]
  wire [3:0] _GEN_457 = 7'h34 == _char_index_1_T_1[6:0] ? 4'h7 : _GEN_456; // @[CharOutput.scala 83:{19,19}]
  wire [3:0] _GEN_458 = 7'h35 == _char_index_1_T_1[6:0] ? 4'h8 : _GEN_457; // @[CharOutput.scala 83:{19,19}]
  wire [3:0] _GEN_459 = 7'h36 == _char_index_1_T_1[6:0] ? 4'h0 : _GEN_458; // @[CharOutput.scala 83:{19,19}]
  wire [3:0] _GEN_460 = 7'h37 == _char_index_1_T_1[6:0] ? 4'h1 : _GEN_459; // @[CharOutput.scala 83:{19,19}]
  wire [3:0] _GEN_461 = 7'h38 == _char_index_1_T_1[6:0] ? 4'h2 : _GEN_460; // @[CharOutput.scala 83:{19,19}]
  wire [3:0] _GEN_462 = 7'h39 == _char_index_1_T_1[6:0] ? 4'h3 : _GEN_461; // @[CharOutput.scala 83:{19,19}]
  wire [3:0] _GEN_463 = 7'h3a == _char_index_1_T_1[6:0] ? 4'h4 : _GEN_462; // @[CharOutput.scala 83:{19,19}]
  wire [3:0] _GEN_464 = 7'h3b == _char_index_1_T_1[6:0] ? 4'h5 : _GEN_463; // @[CharOutput.scala 83:{19,19}]
  wire [3:0] _GEN_465 = 7'h3c == _char_index_1_T_1[6:0] ? 4'h6 : _GEN_464; // @[CharOutput.scala 83:{19,19}]
  wire [3:0] _GEN_466 = 7'h3d == _char_index_1_T_1[6:0] ? 4'h7 : _GEN_465; // @[CharOutput.scala 83:{19,19}]
  wire [3:0] _GEN_467 = 7'h3e == _char_index_1_T_1[6:0] ? 4'h8 : _GEN_466; // @[CharOutput.scala 83:{19,19}]
  wire [3:0] _GEN_468 = 7'h3f == _char_index_1_T_1[6:0] ? 4'h0 : _GEN_467; // @[CharOutput.scala 83:{19,19}]
  wire [3:0] _GEN_469 = 7'h40 == _char_index_1_T_1[6:0] ? 4'h1 : _GEN_468; // @[CharOutput.scala 83:{19,19}]
  wire [3:0] _GEN_470 = 7'h41 == _char_index_1_T_1[6:0] ? 4'h2 : _GEN_469; // @[CharOutput.scala 83:{19,19}]
  wire [3:0] _GEN_471 = 7'h42 == _char_index_1_T_1[6:0] ? 4'h3 : _GEN_470; // @[CharOutput.scala 83:{19,19}]
  wire [3:0] _GEN_472 = 7'h43 == _char_index_1_T_1[6:0] ? 4'h4 : _GEN_471; // @[CharOutput.scala 83:{19,19}]
  wire [3:0] _GEN_473 = 7'h44 == _char_index_1_T_1[6:0] ? 4'h5 : _GEN_472; // @[CharOutput.scala 83:{19,19}]
  wire [3:0] _GEN_474 = 7'h45 == _char_index_1_T_1[6:0] ? 4'h6 : _GEN_473; // @[CharOutput.scala 83:{19,19}]
  wire [3:0] _GEN_475 = 7'h46 == _char_index_1_T_1[6:0] ? 4'h7 : _GEN_474; // @[CharOutput.scala 83:{19,19}]
  wire [3:0] _GEN_476 = 7'h47 == _char_index_1_T_1[6:0] ? 4'h8 : _GEN_475; // @[CharOutput.scala 83:{19,19}]
  wire [3:0] _GEN_477 = 7'h48 == _char_index_1_T_1[6:0] ? 4'h0 : _GEN_476; // @[CharOutput.scala 83:{19,19}]
  wire [3:0] _GEN_478 = 7'h49 == _char_index_1_T_1[6:0] ? 4'h1 : _GEN_477; // @[CharOutput.scala 83:{19,19}]
  wire [3:0] _GEN_479 = 7'h4a == _char_index_1_T_1[6:0] ? 4'h2 : _GEN_478; // @[CharOutput.scala 83:{19,19}]
  wire [3:0] _GEN_480 = 7'h4b == _char_index_1_T_1[6:0] ? 4'h3 : _GEN_479; // @[CharOutput.scala 83:{19,19}]
  wire [3:0] _GEN_481 = 7'h4c == _char_index_1_T_1[6:0] ? 4'h4 : _GEN_480; // @[CharOutput.scala 83:{19,19}]
  wire [3:0] _GEN_482 = 7'h4d == _char_index_1_T_1[6:0] ? 4'h5 : _GEN_481; // @[CharOutput.scala 83:{19,19}]
  wire [3:0] _GEN_483 = 7'h4e == _char_index_1_T_1[6:0] ? 4'h6 : _GEN_482; // @[CharOutput.scala 83:{19,19}]
  wire [3:0] _GEN_484 = 7'h4f == _char_index_1_T_1[6:0] ? 4'h7 : _GEN_483; // @[CharOutput.scala 83:{19,19}]
  wire [3:0] _GEN_485 = 7'h50 == _char_index_1_T_1[6:0] ? 4'h8 : _GEN_484; // @[CharOutput.scala 83:{19,19}]
  wire [3:0] _GEN_486 = 7'h51 == _char_index_1_T_1[6:0] ? 4'h0 : _GEN_485; // @[CharOutput.scala 83:{19,19}]
  wire [3:0] _GEN_487 = 7'h52 == _char_index_1_T_1[6:0] ? 4'h1 : _GEN_486; // @[CharOutput.scala 83:{19,19}]
  wire [3:0] _GEN_488 = 7'h53 == _char_index_1_T_1[6:0] ? 4'h2 : _GEN_487; // @[CharOutput.scala 83:{19,19}]
  wire [3:0] _GEN_489 = 7'h54 == _char_index_1_T_1[6:0] ? 4'h3 : _GEN_488; // @[CharOutput.scala 83:{19,19}]
  wire [3:0] _GEN_490 = 7'h55 == _char_index_1_T_1[6:0] ? 4'h4 : _GEN_489; // @[CharOutput.scala 83:{19,19}]
  wire [3:0] _GEN_491 = 7'h56 == _char_index_1_T_1[6:0] ? 4'h5 : _GEN_490; // @[CharOutput.scala 83:{19,19}]
  wire [3:0] _GEN_492 = 7'h57 == _char_index_1_T_1[6:0] ? 4'h6 : _GEN_491; // @[CharOutput.scala 83:{19,19}]
  wire [3:0] _GEN_493 = 7'h58 == _char_index_1_T_1[6:0] ? 4'h7 : _GEN_492; // @[CharOutput.scala 83:{19,19}]
  wire [3:0] _GEN_494 = 7'h59 == _char_index_1_T_1[6:0] ? 4'h8 : _GEN_493; // @[CharOutput.scala 83:{19,19}]
  wire [3:0] _GEN_495 = 7'h5a == _char_index_1_T_1[6:0] ? 4'h0 : _GEN_494; // @[CharOutput.scala 83:{19,19}]
  wire [3:0] _GEN_496 = 7'h5b == _char_index_1_T_1[6:0] ? 4'h1 : _GEN_495; // @[CharOutput.scala 83:{19,19}]
  wire [3:0] _GEN_497 = 7'h5c == _char_index_1_T_1[6:0] ? 4'h2 : _GEN_496; // @[CharOutput.scala 83:{19,19}]
  wire [3:0] _GEN_498 = 7'h5d == _char_index_1_T_1[6:0] ? 4'h3 : _GEN_497; // @[CharOutput.scala 83:{19,19}]
  wire [3:0] _GEN_499 = 7'h5e == _char_index_1_T_1[6:0] ? 4'h4 : _GEN_498; // @[CharOutput.scala 83:{19,19}]
  wire [3:0] _GEN_500 = 7'h5f == _char_index_1_T_1[6:0] ? 4'h5 : _GEN_499; // @[CharOutput.scala 83:{19,19}]
  wire [3:0] _GEN_501 = 7'h60 == _char_index_1_T_1[6:0] ? 4'h6 : _GEN_500; // @[CharOutput.scala 83:{19,19}]
  wire [3:0] _GEN_502 = 7'h61 == _char_index_1_T_1[6:0] ? 4'h7 : _GEN_501; // @[CharOutput.scala 83:{19,19}]
  wire [3:0] _GEN_503 = 7'h62 == _char_index_1_T_1[6:0] ? 4'h8 : _GEN_502; // @[CharOutput.scala 83:{19,19}]
  wire [3:0] char_index_1 = in_area_h_1 ? _GEN_404 : 4'h0; // @[CharOutput.scala 81:23 82:21 85:21]
  wire [3:0] char_col_1 = in_area_h_1 ? _GEN_503 : 4'h0; // @[CharOutput.scala 81:23 83:19 86:19]
  wire [10:0] _char_row_1_T_1 = io_v_cnt - char_area_ytop_1; // @[CharOutput.scala 89:31]
  wire [10:0] _GEN_506 = in_area_v_1 ? _char_row_1_T_1 : 11'h0; // @[CharOutput.scala 88:23 89:19 91:19]
  wire [10:0] _char_index_2_T_1 = io_h_cnt - io_rect_xleft_2; // @[CharOutput.scala 82:48]
  wire [3:0] _GEN_516 = 7'h9 == _char_index_2_T_1[6:0] ? 4'h1 : 4'h0; // @[CharOutput.scala 82:{21,21}]
  wire [3:0] _GEN_517 = 7'ha == _char_index_2_T_1[6:0] ? 4'h1 : _GEN_516; // @[CharOutput.scala 82:{21,21}]
  wire [3:0] _GEN_518 = 7'hb == _char_index_2_T_1[6:0] ? 4'h1 : _GEN_517; // @[CharOutput.scala 82:{21,21}]
  wire [3:0] _GEN_519 = 7'hc == _char_index_2_T_1[6:0] ? 4'h1 : _GEN_518; // @[CharOutput.scala 82:{21,21}]
  wire [3:0] _GEN_520 = 7'hd == _char_index_2_T_1[6:0] ? 4'h1 : _GEN_519; // @[CharOutput.scala 82:{21,21}]
  wire [3:0] _GEN_521 = 7'he == _char_index_2_T_1[6:0] ? 4'h1 : _GEN_520; // @[CharOutput.scala 82:{21,21}]
  wire [3:0] _GEN_522 = 7'hf == _char_index_2_T_1[6:0] ? 4'h1 : _GEN_521; // @[CharOutput.scala 82:{21,21}]
  wire [3:0] _GEN_523 = 7'h10 == _char_index_2_T_1[6:0] ? 4'h1 : _GEN_522; // @[CharOutput.scala 82:{21,21}]
  wire [3:0] _GEN_524 = 7'h11 == _char_index_2_T_1[6:0] ? 4'h1 : _GEN_523; // @[CharOutput.scala 82:{21,21}]
  wire [3:0] _GEN_525 = 7'h12 == _char_index_2_T_1[6:0] ? 4'h2 : _GEN_524; // @[CharOutput.scala 82:{21,21}]
  wire [3:0] _GEN_526 = 7'h13 == _char_index_2_T_1[6:0] ? 4'h2 : _GEN_525; // @[CharOutput.scala 82:{21,21}]
  wire [3:0] _GEN_527 = 7'h14 == _char_index_2_T_1[6:0] ? 4'h2 : _GEN_526; // @[CharOutput.scala 82:{21,21}]
  wire [3:0] _GEN_528 = 7'h15 == _char_index_2_T_1[6:0] ? 4'h2 : _GEN_527; // @[CharOutput.scala 82:{21,21}]
  wire [3:0] _GEN_529 = 7'h16 == _char_index_2_T_1[6:0] ? 4'h2 : _GEN_528; // @[CharOutput.scala 82:{21,21}]
  wire [3:0] _GEN_530 = 7'h17 == _char_index_2_T_1[6:0] ? 4'h2 : _GEN_529; // @[CharOutput.scala 82:{21,21}]
  wire [3:0] _GEN_531 = 7'h18 == _char_index_2_T_1[6:0] ? 4'h2 : _GEN_530; // @[CharOutput.scala 82:{21,21}]
  wire [3:0] _GEN_532 = 7'h19 == _char_index_2_T_1[6:0] ? 4'h2 : _GEN_531; // @[CharOutput.scala 82:{21,21}]
  wire [3:0] _GEN_533 = 7'h1a == _char_index_2_T_1[6:0] ? 4'h2 : _GEN_532; // @[CharOutput.scala 82:{21,21}]
  wire [3:0] _GEN_534 = 7'h1b == _char_index_2_T_1[6:0] ? 4'h3 : _GEN_533; // @[CharOutput.scala 82:{21,21}]
  wire [3:0] _GEN_535 = 7'h1c == _char_index_2_T_1[6:0] ? 4'h3 : _GEN_534; // @[CharOutput.scala 82:{21,21}]
  wire [3:0] _GEN_536 = 7'h1d == _char_index_2_T_1[6:0] ? 4'h3 : _GEN_535; // @[CharOutput.scala 82:{21,21}]
  wire [3:0] _GEN_537 = 7'h1e == _char_index_2_T_1[6:0] ? 4'h3 : _GEN_536; // @[CharOutput.scala 82:{21,21}]
  wire [3:0] _GEN_538 = 7'h1f == _char_index_2_T_1[6:0] ? 4'h3 : _GEN_537; // @[CharOutput.scala 82:{21,21}]
  wire [3:0] _GEN_539 = 7'h20 == _char_index_2_T_1[6:0] ? 4'h3 : _GEN_538; // @[CharOutput.scala 82:{21,21}]
  wire [3:0] _GEN_540 = 7'h21 == _char_index_2_T_1[6:0] ? 4'h3 : _GEN_539; // @[CharOutput.scala 82:{21,21}]
  wire [3:0] _GEN_541 = 7'h22 == _char_index_2_T_1[6:0] ? 4'h3 : _GEN_540; // @[CharOutput.scala 82:{21,21}]
  wire [3:0] _GEN_542 = 7'h23 == _char_index_2_T_1[6:0] ? 4'h3 : _GEN_541; // @[CharOutput.scala 82:{21,21}]
  wire [3:0] _GEN_543 = 7'h24 == _char_index_2_T_1[6:0] ? 4'h4 : _GEN_542; // @[CharOutput.scala 82:{21,21}]
  wire [3:0] _GEN_544 = 7'h25 == _char_index_2_T_1[6:0] ? 4'h4 : _GEN_543; // @[CharOutput.scala 82:{21,21}]
  wire [3:0] _GEN_545 = 7'h26 == _char_index_2_T_1[6:0] ? 4'h4 : _GEN_544; // @[CharOutput.scala 82:{21,21}]
  wire [3:0] _GEN_546 = 7'h27 == _char_index_2_T_1[6:0] ? 4'h4 : _GEN_545; // @[CharOutput.scala 82:{21,21}]
  wire [3:0] _GEN_547 = 7'h28 == _char_index_2_T_1[6:0] ? 4'h4 : _GEN_546; // @[CharOutput.scala 82:{21,21}]
  wire [3:0] _GEN_548 = 7'h29 == _char_index_2_T_1[6:0] ? 4'h4 : _GEN_547; // @[CharOutput.scala 82:{21,21}]
  wire [3:0] _GEN_549 = 7'h2a == _char_index_2_T_1[6:0] ? 4'h4 : _GEN_548; // @[CharOutput.scala 82:{21,21}]
  wire [3:0] _GEN_550 = 7'h2b == _char_index_2_T_1[6:0] ? 4'h4 : _GEN_549; // @[CharOutput.scala 82:{21,21}]
  wire [3:0] _GEN_551 = 7'h2c == _char_index_2_T_1[6:0] ? 4'h4 : _GEN_550; // @[CharOutput.scala 82:{21,21}]
  wire [3:0] _GEN_552 = 7'h2d == _char_index_2_T_1[6:0] ? 4'h5 : _GEN_551; // @[CharOutput.scala 82:{21,21}]
  wire [3:0] _GEN_553 = 7'h2e == _char_index_2_T_1[6:0] ? 4'h5 : _GEN_552; // @[CharOutput.scala 82:{21,21}]
  wire [3:0] _GEN_554 = 7'h2f == _char_index_2_T_1[6:0] ? 4'h5 : _GEN_553; // @[CharOutput.scala 82:{21,21}]
  wire [3:0] _GEN_555 = 7'h30 == _char_index_2_T_1[6:0] ? 4'h5 : _GEN_554; // @[CharOutput.scala 82:{21,21}]
  wire [3:0] _GEN_556 = 7'h31 == _char_index_2_T_1[6:0] ? 4'h5 : _GEN_555; // @[CharOutput.scala 82:{21,21}]
  wire [3:0] _GEN_557 = 7'h32 == _char_index_2_T_1[6:0] ? 4'h5 : _GEN_556; // @[CharOutput.scala 82:{21,21}]
  wire [3:0] _GEN_558 = 7'h33 == _char_index_2_T_1[6:0] ? 4'h5 : _GEN_557; // @[CharOutput.scala 82:{21,21}]
  wire [3:0] _GEN_559 = 7'h34 == _char_index_2_T_1[6:0] ? 4'h5 : _GEN_558; // @[CharOutput.scala 82:{21,21}]
  wire [3:0] _GEN_560 = 7'h35 == _char_index_2_T_1[6:0] ? 4'h5 : _GEN_559; // @[CharOutput.scala 82:{21,21}]
  wire [3:0] _GEN_561 = 7'h36 == _char_index_2_T_1[6:0] ? 4'h6 : _GEN_560; // @[CharOutput.scala 82:{21,21}]
  wire [3:0] _GEN_562 = 7'h37 == _char_index_2_T_1[6:0] ? 4'h6 : _GEN_561; // @[CharOutput.scala 82:{21,21}]
  wire [3:0] _GEN_563 = 7'h38 == _char_index_2_T_1[6:0] ? 4'h6 : _GEN_562; // @[CharOutput.scala 82:{21,21}]
  wire [3:0] _GEN_564 = 7'h39 == _char_index_2_T_1[6:0] ? 4'h6 : _GEN_563; // @[CharOutput.scala 82:{21,21}]
  wire [3:0] _GEN_565 = 7'h3a == _char_index_2_T_1[6:0] ? 4'h6 : _GEN_564; // @[CharOutput.scala 82:{21,21}]
  wire [3:0] _GEN_566 = 7'h3b == _char_index_2_T_1[6:0] ? 4'h6 : _GEN_565; // @[CharOutput.scala 82:{21,21}]
  wire [3:0] _GEN_567 = 7'h3c == _char_index_2_T_1[6:0] ? 4'h6 : _GEN_566; // @[CharOutput.scala 82:{21,21}]
  wire [3:0] _GEN_568 = 7'h3d == _char_index_2_T_1[6:0] ? 4'h6 : _GEN_567; // @[CharOutput.scala 82:{21,21}]
  wire [3:0] _GEN_569 = 7'h3e == _char_index_2_T_1[6:0] ? 4'h6 : _GEN_568; // @[CharOutput.scala 82:{21,21}]
  wire [3:0] _GEN_570 = 7'h3f == _char_index_2_T_1[6:0] ? 4'h7 : _GEN_569; // @[CharOutput.scala 82:{21,21}]
  wire [3:0] _GEN_571 = 7'h40 == _char_index_2_T_1[6:0] ? 4'h7 : _GEN_570; // @[CharOutput.scala 82:{21,21}]
  wire [3:0] _GEN_572 = 7'h41 == _char_index_2_T_1[6:0] ? 4'h7 : _GEN_571; // @[CharOutput.scala 82:{21,21}]
  wire [3:0] _GEN_573 = 7'h42 == _char_index_2_T_1[6:0] ? 4'h7 : _GEN_572; // @[CharOutput.scala 82:{21,21}]
  wire [3:0] _GEN_574 = 7'h43 == _char_index_2_T_1[6:0] ? 4'h7 : _GEN_573; // @[CharOutput.scala 82:{21,21}]
  wire [3:0] _GEN_575 = 7'h44 == _char_index_2_T_1[6:0] ? 4'h7 : _GEN_574; // @[CharOutput.scala 82:{21,21}]
  wire [3:0] _GEN_576 = 7'h45 == _char_index_2_T_1[6:0] ? 4'h7 : _GEN_575; // @[CharOutput.scala 82:{21,21}]
  wire [3:0] _GEN_577 = 7'h46 == _char_index_2_T_1[6:0] ? 4'h7 : _GEN_576; // @[CharOutput.scala 82:{21,21}]
  wire [3:0] _GEN_578 = 7'h47 == _char_index_2_T_1[6:0] ? 4'h7 : _GEN_577; // @[CharOutput.scala 82:{21,21}]
  wire [3:0] _GEN_579 = 7'h48 == _char_index_2_T_1[6:0] ? 4'h8 : _GEN_578; // @[CharOutput.scala 82:{21,21}]
  wire [3:0] _GEN_580 = 7'h49 == _char_index_2_T_1[6:0] ? 4'h8 : _GEN_579; // @[CharOutput.scala 82:{21,21}]
  wire [3:0] _GEN_581 = 7'h4a == _char_index_2_T_1[6:0] ? 4'h8 : _GEN_580; // @[CharOutput.scala 82:{21,21}]
  wire [3:0] _GEN_582 = 7'h4b == _char_index_2_T_1[6:0] ? 4'h8 : _GEN_581; // @[CharOutput.scala 82:{21,21}]
  wire [3:0] _GEN_583 = 7'h4c == _char_index_2_T_1[6:0] ? 4'h8 : _GEN_582; // @[CharOutput.scala 82:{21,21}]
  wire [3:0] _GEN_584 = 7'h4d == _char_index_2_T_1[6:0] ? 4'h8 : _GEN_583; // @[CharOutput.scala 82:{21,21}]
  wire [3:0] _GEN_585 = 7'h4e == _char_index_2_T_1[6:0] ? 4'h8 : _GEN_584; // @[CharOutput.scala 82:{21,21}]
  wire [3:0] _GEN_586 = 7'h4f == _char_index_2_T_1[6:0] ? 4'h8 : _GEN_585; // @[CharOutput.scala 82:{21,21}]
  wire [3:0] _GEN_587 = 7'h50 == _char_index_2_T_1[6:0] ? 4'h8 : _GEN_586; // @[CharOutput.scala 82:{21,21}]
  wire [3:0] _GEN_588 = 7'h51 == _char_index_2_T_1[6:0] ? 4'h9 : _GEN_587; // @[CharOutput.scala 82:{21,21}]
  wire [3:0] _GEN_589 = 7'h52 == _char_index_2_T_1[6:0] ? 4'h9 : _GEN_588; // @[CharOutput.scala 82:{21,21}]
  wire [3:0] _GEN_590 = 7'h53 == _char_index_2_T_1[6:0] ? 4'h9 : _GEN_589; // @[CharOutput.scala 82:{21,21}]
  wire [3:0] _GEN_591 = 7'h54 == _char_index_2_T_1[6:0] ? 4'h9 : _GEN_590; // @[CharOutput.scala 82:{21,21}]
  wire [3:0] _GEN_592 = 7'h55 == _char_index_2_T_1[6:0] ? 4'h9 : _GEN_591; // @[CharOutput.scala 82:{21,21}]
  wire [3:0] _GEN_593 = 7'h56 == _char_index_2_T_1[6:0] ? 4'h9 : _GEN_592; // @[CharOutput.scala 82:{21,21}]
  wire [3:0] _GEN_594 = 7'h57 == _char_index_2_T_1[6:0] ? 4'h9 : _GEN_593; // @[CharOutput.scala 82:{21,21}]
  wire [3:0] _GEN_595 = 7'h58 == _char_index_2_T_1[6:0] ? 4'h9 : _GEN_594; // @[CharOutput.scala 82:{21,21}]
  wire [3:0] _GEN_596 = 7'h59 == _char_index_2_T_1[6:0] ? 4'h9 : _GEN_595; // @[CharOutput.scala 82:{21,21}]
  wire [3:0] _GEN_597 = 7'h5a == _char_index_2_T_1[6:0] ? 4'ha : _GEN_596; // @[CharOutput.scala 82:{21,21}]
  wire [3:0] _GEN_598 = 7'h5b == _char_index_2_T_1[6:0] ? 4'ha : _GEN_597; // @[CharOutput.scala 82:{21,21}]
  wire [3:0] _GEN_599 = 7'h5c == _char_index_2_T_1[6:0] ? 4'ha : _GEN_598; // @[CharOutput.scala 82:{21,21}]
  wire [3:0] _GEN_600 = 7'h5d == _char_index_2_T_1[6:0] ? 4'ha : _GEN_599; // @[CharOutput.scala 82:{21,21}]
  wire [3:0] _GEN_601 = 7'h5e == _char_index_2_T_1[6:0] ? 4'ha : _GEN_600; // @[CharOutput.scala 82:{21,21}]
  wire [3:0] _GEN_602 = 7'h5f == _char_index_2_T_1[6:0] ? 4'ha : _GEN_601; // @[CharOutput.scala 82:{21,21}]
  wire [3:0] _GEN_603 = 7'h60 == _char_index_2_T_1[6:0] ? 4'ha : _GEN_602; // @[CharOutput.scala 82:{21,21}]
  wire [3:0] _GEN_604 = 7'h61 == _char_index_2_T_1[6:0] ? 4'ha : _GEN_603; // @[CharOutput.scala 82:{21,21}]
  wire [3:0] _GEN_605 = 7'h62 == _char_index_2_T_1[6:0] ? 4'ha : _GEN_604; // @[CharOutput.scala 82:{21,21}]
  wire [3:0] _GEN_607 = 7'h1 == _char_index_2_T_1[6:0] ? 4'h1 : 4'h0; // @[CharOutput.scala 83:{19,19}]
  wire [3:0] _GEN_608 = 7'h2 == _char_index_2_T_1[6:0] ? 4'h2 : _GEN_607; // @[CharOutput.scala 83:{19,19}]
  wire [3:0] _GEN_609 = 7'h3 == _char_index_2_T_1[6:0] ? 4'h3 : _GEN_608; // @[CharOutput.scala 83:{19,19}]
  wire [3:0] _GEN_610 = 7'h4 == _char_index_2_T_1[6:0] ? 4'h4 : _GEN_609; // @[CharOutput.scala 83:{19,19}]
  wire [3:0] _GEN_611 = 7'h5 == _char_index_2_T_1[6:0] ? 4'h5 : _GEN_610; // @[CharOutput.scala 83:{19,19}]
  wire [3:0] _GEN_612 = 7'h6 == _char_index_2_T_1[6:0] ? 4'h6 : _GEN_611; // @[CharOutput.scala 83:{19,19}]
  wire [3:0] _GEN_613 = 7'h7 == _char_index_2_T_1[6:0] ? 4'h7 : _GEN_612; // @[CharOutput.scala 83:{19,19}]
  wire [3:0] _GEN_614 = 7'h8 == _char_index_2_T_1[6:0] ? 4'h8 : _GEN_613; // @[CharOutput.scala 83:{19,19}]
  wire [3:0] _GEN_615 = 7'h9 == _char_index_2_T_1[6:0] ? 4'h0 : _GEN_614; // @[CharOutput.scala 83:{19,19}]
  wire [3:0] _GEN_616 = 7'ha == _char_index_2_T_1[6:0] ? 4'h1 : _GEN_615; // @[CharOutput.scala 83:{19,19}]
  wire [3:0] _GEN_617 = 7'hb == _char_index_2_T_1[6:0] ? 4'h2 : _GEN_616; // @[CharOutput.scala 83:{19,19}]
  wire [3:0] _GEN_618 = 7'hc == _char_index_2_T_1[6:0] ? 4'h3 : _GEN_617; // @[CharOutput.scala 83:{19,19}]
  wire [3:0] _GEN_619 = 7'hd == _char_index_2_T_1[6:0] ? 4'h4 : _GEN_618; // @[CharOutput.scala 83:{19,19}]
  wire [3:0] _GEN_620 = 7'he == _char_index_2_T_1[6:0] ? 4'h5 : _GEN_619; // @[CharOutput.scala 83:{19,19}]
  wire [3:0] _GEN_621 = 7'hf == _char_index_2_T_1[6:0] ? 4'h6 : _GEN_620; // @[CharOutput.scala 83:{19,19}]
  wire [3:0] _GEN_622 = 7'h10 == _char_index_2_T_1[6:0] ? 4'h7 : _GEN_621; // @[CharOutput.scala 83:{19,19}]
  wire [3:0] _GEN_623 = 7'h11 == _char_index_2_T_1[6:0] ? 4'h8 : _GEN_622; // @[CharOutput.scala 83:{19,19}]
  wire [3:0] _GEN_624 = 7'h12 == _char_index_2_T_1[6:0] ? 4'h0 : _GEN_623; // @[CharOutput.scala 83:{19,19}]
  wire [3:0] _GEN_625 = 7'h13 == _char_index_2_T_1[6:0] ? 4'h1 : _GEN_624; // @[CharOutput.scala 83:{19,19}]
  wire [3:0] _GEN_626 = 7'h14 == _char_index_2_T_1[6:0] ? 4'h2 : _GEN_625; // @[CharOutput.scala 83:{19,19}]
  wire [3:0] _GEN_627 = 7'h15 == _char_index_2_T_1[6:0] ? 4'h3 : _GEN_626; // @[CharOutput.scala 83:{19,19}]
  wire [3:0] _GEN_628 = 7'h16 == _char_index_2_T_1[6:0] ? 4'h4 : _GEN_627; // @[CharOutput.scala 83:{19,19}]
  wire [3:0] _GEN_629 = 7'h17 == _char_index_2_T_1[6:0] ? 4'h5 : _GEN_628; // @[CharOutput.scala 83:{19,19}]
  wire [3:0] _GEN_630 = 7'h18 == _char_index_2_T_1[6:0] ? 4'h6 : _GEN_629; // @[CharOutput.scala 83:{19,19}]
  wire [3:0] _GEN_631 = 7'h19 == _char_index_2_T_1[6:0] ? 4'h7 : _GEN_630; // @[CharOutput.scala 83:{19,19}]
  wire [3:0] _GEN_632 = 7'h1a == _char_index_2_T_1[6:0] ? 4'h8 : _GEN_631; // @[CharOutput.scala 83:{19,19}]
  wire [3:0] _GEN_633 = 7'h1b == _char_index_2_T_1[6:0] ? 4'h0 : _GEN_632; // @[CharOutput.scala 83:{19,19}]
  wire [3:0] _GEN_634 = 7'h1c == _char_index_2_T_1[6:0] ? 4'h1 : _GEN_633; // @[CharOutput.scala 83:{19,19}]
  wire [3:0] _GEN_635 = 7'h1d == _char_index_2_T_1[6:0] ? 4'h2 : _GEN_634; // @[CharOutput.scala 83:{19,19}]
  wire [3:0] _GEN_636 = 7'h1e == _char_index_2_T_1[6:0] ? 4'h3 : _GEN_635; // @[CharOutput.scala 83:{19,19}]
  wire [3:0] _GEN_637 = 7'h1f == _char_index_2_T_1[6:0] ? 4'h4 : _GEN_636; // @[CharOutput.scala 83:{19,19}]
  wire [3:0] _GEN_638 = 7'h20 == _char_index_2_T_1[6:0] ? 4'h5 : _GEN_637; // @[CharOutput.scala 83:{19,19}]
  wire [3:0] _GEN_639 = 7'h21 == _char_index_2_T_1[6:0] ? 4'h6 : _GEN_638; // @[CharOutput.scala 83:{19,19}]
  wire [3:0] _GEN_640 = 7'h22 == _char_index_2_T_1[6:0] ? 4'h7 : _GEN_639; // @[CharOutput.scala 83:{19,19}]
  wire [3:0] _GEN_641 = 7'h23 == _char_index_2_T_1[6:0] ? 4'h8 : _GEN_640; // @[CharOutput.scala 83:{19,19}]
  wire [3:0] _GEN_642 = 7'h24 == _char_index_2_T_1[6:0] ? 4'h0 : _GEN_641; // @[CharOutput.scala 83:{19,19}]
  wire [3:0] _GEN_643 = 7'h25 == _char_index_2_T_1[6:0] ? 4'h1 : _GEN_642; // @[CharOutput.scala 83:{19,19}]
  wire [3:0] _GEN_644 = 7'h26 == _char_index_2_T_1[6:0] ? 4'h2 : _GEN_643; // @[CharOutput.scala 83:{19,19}]
  wire [3:0] _GEN_645 = 7'h27 == _char_index_2_T_1[6:0] ? 4'h3 : _GEN_644; // @[CharOutput.scala 83:{19,19}]
  wire [3:0] _GEN_646 = 7'h28 == _char_index_2_T_1[6:0] ? 4'h4 : _GEN_645; // @[CharOutput.scala 83:{19,19}]
  wire [3:0] _GEN_647 = 7'h29 == _char_index_2_T_1[6:0] ? 4'h5 : _GEN_646; // @[CharOutput.scala 83:{19,19}]
  wire [3:0] _GEN_648 = 7'h2a == _char_index_2_T_1[6:0] ? 4'h6 : _GEN_647; // @[CharOutput.scala 83:{19,19}]
  wire [3:0] _GEN_649 = 7'h2b == _char_index_2_T_1[6:0] ? 4'h7 : _GEN_648; // @[CharOutput.scala 83:{19,19}]
  wire [3:0] _GEN_650 = 7'h2c == _char_index_2_T_1[6:0] ? 4'h8 : _GEN_649; // @[CharOutput.scala 83:{19,19}]
  wire [3:0] _GEN_651 = 7'h2d == _char_index_2_T_1[6:0] ? 4'h0 : _GEN_650; // @[CharOutput.scala 83:{19,19}]
  wire [3:0] _GEN_652 = 7'h2e == _char_index_2_T_1[6:0] ? 4'h1 : _GEN_651; // @[CharOutput.scala 83:{19,19}]
  wire [3:0] _GEN_653 = 7'h2f == _char_index_2_T_1[6:0] ? 4'h2 : _GEN_652; // @[CharOutput.scala 83:{19,19}]
  wire [3:0] _GEN_654 = 7'h30 == _char_index_2_T_1[6:0] ? 4'h3 : _GEN_653; // @[CharOutput.scala 83:{19,19}]
  wire [3:0] _GEN_655 = 7'h31 == _char_index_2_T_1[6:0] ? 4'h4 : _GEN_654; // @[CharOutput.scala 83:{19,19}]
  wire [3:0] _GEN_656 = 7'h32 == _char_index_2_T_1[6:0] ? 4'h5 : _GEN_655; // @[CharOutput.scala 83:{19,19}]
  wire [3:0] _GEN_657 = 7'h33 == _char_index_2_T_1[6:0] ? 4'h6 : _GEN_656; // @[CharOutput.scala 83:{19,19}]
  wire [3:0] _GEN_658 = 7'h34 == _char_index_2_T_1[6:0] ? 4'h7 : _GEN_657; // @[CharOutput.scala 83:{19,19}]
  wire [3:0] _GEN_659 = 7'h35 == _char_index_2_T_1[6:0] ? 4'h8 : _GEN_658; // @[CharOutput.scala 83:{19,19}]
  wire [3:0] _GEN_660 = 7'h36 == _char_index_2_T_1[6:0] ? 4'h0 : _GEN_659; // @[CharOutput.scala 83:{19,19}]
  wire [3:0] _GEN_661 = 7'h37 == _char_index_2_T_1[6:0] ? 4'h1 : _GEN_660; // @[CharOutput.scala 83:{19,19}]
  wire [3:0] _GEN_662 = 7'h38 == _char_index_2_T_1[6:0] ? 4'h2 : _GEN_661; // @[CharOutput.scala 83:{19,19}]
  wire [3:0] _GEN_663 = 7'h39 == _char_index_2_T_1[6:0] ? 4'h3 : _GEN_662; // @[CharOutput.scala 83:{19,19}]
  wire [3:0] _GEN_664 = 7'h3a == _char_index_2_T_1[6:0] ? 4'h4 : _GEN_663; // @[CharOutput.scala 83:{19,19}]
  wire [3:0] _GEN_665 = 7'h3b == _char_index_2_T_1[6:0] ? 4'h5 : _GEN_664; // @[CharOutput.scala 83:{19,19}]
  wire [3:0] _GEN_666 = 7'h3c == _char_index_2_T_1[6:0] ? 4'h6 : _GEN_665; // @[CharOutput.scala 83:{19,19}]
  wire [3:0] _GEN_667 = 7'h3d == _char_index_2_T_1[6:0] ? 4'h7 : _GEN_666; // @[CharOutput.scala 83:{19,19}]
  wire [3:0] _GEN_668 = 7'h3e == _char_index_2_T_1[6:0] ? 4'h8 : _GEN_667; // @[CharOutput.scala 83:{19,19}]
  wire [3:0] _GEN_669 = 7'h3f == _char_index_2_T_1[6:0] ? 4'h0 : _GEN_668; // @[CharOutput.scala 83:{19,19}]
  wire [3:0] _GEN_670 = 7'h40 == _char_index_2_T_1[6:0] ? 4'h1 : _GEN_669; // @[CharOutput.scala 83:{19,19}]
  wire [3:0] _GEN_671 = 7'h41 == _char_index_2_T_1[6:0] ? 4'h2 : _GEN_670; // @[CharOutput.scala 83:{19,19}]
  wire [3:0] _GEN_672 = 7'h42 == _char_index_2_T_1[6:0] ? 4'h3 : _GEN_671; // @[CharOutput.scala 83:{19,19}]
  wire [3:0] _GEN_673 = 7'h43 == _char_index_2_T_1[6:0] ? 4'h4 : _GEN_672; // @[CharOutput.scala 83:{19,19}]
  wire [3:0] _GEN_674 = 7'h44 == _char_index_2_T_1[6:0] ? 4'h5 : _GEN_673; // @[CharOutput.scala 83:{19,19}]
  wire [3:0] _GEN_675 = 7'h45 == _char_index_2_T_1[6:0] ? 4'h6 : _GEN_674; // @[CharOutput.scala 83:{19,19}]
  wire [3:0] _GEN_676 = 7'h46 == _char_index_2_T_1[6:0] ? 4'h7 : _GEN_675; // @[CharOutput.scala 83:{19,19}]
  wire [3:0] _GEN_677 = 7'h47 == _char_index_2_T_1[6:0] ? 4'h8 : _GEN_676; // @[CharOutput.scala 83:{19,19}]
  wire [3:0] _GEN_678 = 7'h48 == _char_index_2_T_1[6:0] ? 4'h0 : _GEN_677; // @[CharOutput.scala 83:{19,19}]
  wire [3:0] _GEN_679 = 7'h49 == _char_index_2_T_1[6:0] ? 4'h1 : _GEN_678; // @[CharOutput.scala 83:{19,19}]
  wire [3:0] _GEN_680 = 7'h4a == _char_index_2_T_1[6:0] ? 4'h2 : _GEN_679; // @[CharOutput.scala 83:{19,19}]
  wire [3:0] _GEN_681 = 7'h4b == _char_index_2_T_1[6:0] ? 4'h3 : _GEN_680; // @[CharOutput.scala 83:{19,19}]
  wire [3:0] _GEN_682 = 7'h4c == _char_index_2_T_1[6:0] ? 4'h4 : _GEN_681; // @[CharOutput.scala 83:{19,19}]
  wire [3:0] _GEN_683 = 7'h4d == _char_index_2_T_1[6:0] ? 4'h5 : _GEN_682; // @[CharOutput.scala 83:{19,19}]
  wire [3:0] _GEN_684 = 7'h4e == _char_index_2_T_1[6:0] ? 4'h6 : _GEN_683; // @[CharOutput.scala 83:{19,19}]
  wire [3:0] _GEN_685 = 7'h4f == _char_index_2_T_1[6:0] ? 4'h7 : _GEN_684; // @[CharOutput.scala 83:{19,19}]
  wire [3:0] _GEN_686 = 7'h50 == _char_index_2_T_1[6:0] ? 4'h8 : _GEN_685; // @[CharOutput.scala 83:{19,19}]
  wire [3:0] _GEN_687 = 7'h51 == _char_index_2_T_1[6:0] ? 4'h0 : _GEN_686; // @[CharOutput.scala 83:{19,19}]
  wire [3:0] _GEN_688 = 7'h52 == _char_index_2_T_1[6:0] ? 4'h1 : _GEN_687; // @[CharOutput.scala 83:{19,19}]
  wire [3:0] _GEN_689 = 7'h53 == _char_index_2_T_1[6:0] ? 4'h2 : _GEN_688; // @[CharOutput.scala 83:{19,19}]
  wire [3:0] _GEN_690 = 7'h54 == _char_index_2_T_1[6:0] ? 4'h3 : _GEN_689; // @[CharOutput.scala 83:{19,19}]
  wire [3:0] _GEN_691 = 7'h55 == _char_index_2_T_1[6:0] ? 4'h4 : _GEN_690; // @[CharOutput.scala 83:{19,19}]
  wire [3:0] _GEN_692 = 7'h56 == _char_index_2_T_1[6:0] ? 4'h5 : _GEN_691; // @[CharOutput.scala 83:{19,19}]
  wire [3:0] _GEN_693 = 7'h57 == _char_index_2_T_1[6:0] ? 4'h6 : _GEN_692; // @[CharOutput.scala 83:{19,19}]
  wire [3:0] _GEN_694 = 7'h58 == _char_index_2_T_1[6:0] ? 4'h7 : _GEN_693; // @[CharOutput.scala 83:{19,19}]
  wire [3:0] _GEN_695 = 7'h59 == _char_index_2_T_1[6:0] ? 4'h8 : _GEN_694; // @[CharOutput.scala 83:{19,19}]
  wire [3:0] _GEN_696 = 7'h5a == _char_index_2_T_1[6:0] ? 4'h0 : _GEN_695; // @[CharOutput.scala 83:{19,19}]
  wire [3:0] _GEN_697 = 7'h5b == _char_index_2_T_1[6:0] ? 4'h1 : _GEN_696; // @[CharOutput.scala 83:{19,19}]
  wire [3:0] _GEN_698 = 7'h5c == _char_index_2_T_1[6:0] ? 4'h2 : _GEN_697; // @[CharOutput.scala 83:{19,19}]
  wire [3:0] _GEN_699 = 7'h5d == _char_index_2_T_1[6:0] ? 4'h3 : _GEN_698; // @[CharOutput.scala 83:{19,19}]
  wire [3:0] _GEN_700 = 7'h5e == _char_index_2_T_1[6:0] ? 4'h4 : _GEN_699; // @[CharOutput.scala 83:{19,19}]
  wire [3:0] _GEN_701 = 7'h5f == _char_index_2_T_1[6:0] ? 4'h5 : _GEN_700; // @[CharOutput.scala 83:{19,19}]
  wire [3:0] _GEN_702 = 7'h60 == _char_index_2_T_1[6:0] ? 4'h6 : _GEN_701; // @[CharOutput.scala 83:{19,19}]
  wire [3:0] _GEN_703 = 7'h61 == _char_index_2_T_1[6:0] ? 4'h7 : _GEN_702; // @[CharOutput.scala 83:{19,19}]
  wire [3:0] _GEN_704 = 7'h62 == _char_index_2_T_1[6:0] ? 4'h8 : _GEN_703; // @[CharOutput.scala 83:{19,19}]
  wire [3:0] char_index_2 = in_area_h_2 ? _GEN_605 : 4'h0; // @[CharOutput.scala 81:23 82:21 85:21]
  wire [3:0] char_col_2 = in_area_h_2 ? _GEN_704 : 4'h0; // @[CharOutput.scala 81:23 83:19 86:19]
  wire [10:0] _char_row_2_T_1 = io_v_cnt - char_area_ytop_2; // @[CharOutput.scala 89:31]
  wire [10:0] _GEN_707 = in_area_v_2 ? _char_row_2_T_1 : 11'h0; // @[CharOutput.scala 88:23 89:19 91:19]
  wire [10:0] _char_index_3_T_1 = io_h_cnt - io_rect_xleft_3; // @[CharOutput.scala 82:48]
  wire [3:0] _GEN_717 = 7'h9 == _char_index_3_T_1[6:0] ? 4'h1 : 4'h0; // @[CharOutput.scala 82:{21,21}]
  wire [3:0] _GEN_718 = 7'ha == _char_index_3_T_1[6:0] ? 4'h1 : _GEN_717; // @[CharOutput.scala 82:{21,21}]
  wire [3:0] _GEN_719 = 7'hb == _char_index_3_T_1[6:0] ? 4'h1 : _GEN_718; // @[CharOutput.scala 82:{21,21}]
  wire [3:0] _GEN_720 = 7'hc == _char_index_3_T_1[6:0] ? 4'h1 : _GEN_719; // @[CharOutput.scala 82:{21,21}]
  wire [3:0] _GEN_721 = 7'hd == _char_index_3_T_1[6:0] ? 4'h1 : _GEN_720; // @[CharOutput.scala 82:{21,21}]
  wire [3:0] _GEN_722 = 7'he == _char_index_3_T_1[6:0] ? 4'h1 : _GEN_721; // @[CharOutput.scala 82:{21,21}]
  wire [3:0] _GEN_723 = 7'hf == _char_index_3_T_1[6:0] ? 4'h1 : _GEN_722; // @[CharOutput.scala 82:{21,21}]
  wire [3:0] _GEN_724 = 7'h10 == _char_index_3_T_1[6:0] ? 4'h1 : _GEN_723; // @[CharOutput.scala 82:{21,21}]
  wire [3:0] _GEN_725 = 7'h11 == _char_index_3_T_1[6:0] ? 4'h1 : _GEN_724; // @[CharOutput.scala 82:{21,21}]
  wire [3:0] _GEN_726 = 7'h12 == _char_index_3_T_1[6:0] ? 4'h2 : _GEN_725; // @[CharOutput.scala 82:{21,21}]
  wire [3:0] _GEN_727 = 7'h13 == _char_index_3_T_1[6:0] ? 4'h2 : _GEN_726; // @[CharOutput.scala 82:{21,21}]
  wire [3:0] _GEN_728 = 7'h14 == _char_index_3_T_1[6:0] ? 4'h2 : _GEN_727; // @[CharOutput.scala 82:{21,21}]
  wire [3:0] _GEN_729 = 7'h15 == _char_index_3_T_1[6:0] ? 4'h2 : _GEN_728; // @[CharOutput.scala 82:{21,21}]
  wire [3:0] _GEN_730 = 7'h16 == _char_index_3_T_1[6:0] ? 4'h2 : _GEN_729; // @[CharOutput.scala 82:{21,21}]
  wire [3:0] _GEN_731 = 7'h17 == _char_index_3_T_1[6:0] ? 4'h2 : _GEN_730; // @[CharOutput.scala 82:{21,21}]
  wire [3:0] _GEN_732 = 7'h18 == _char_index_3_T_1[6:0] ? 4'h2 : _GEN_731; // @[CharOutput.scala 82:{21,21}]
  wire [3:0] _GEN_733 = 7'h19 == _char_index_3_T_1[6:0] ? 4'h2 : _GEN_732; // @[CharOutput.scala 82:{21,21}]
  wire [3:0] _GEN_734 = 7'h1a == _char_index_3_T_1[6:0] ? 4'h2 : _GEN_733; // @[CharOutput.scala 82:{21,21}]
  wire [3:0] _GEN_735 = 7'h1b == _char_index_3_T_1[6:0] ? 4'h3 : _GEN_734; // @[CharOutput.scala 82:{21,21}]
  wire [3:0] _GEN_736 = 7'h1c == _char_index_3_T_1[6:0] ? 4'h3 : _GEN_735; // @[CharOutput.scala 82:{21,21}]
  wire [3:0] _GEN_737 = 7'h1d == _char_index_3_T_1[6:0] ? 4'h3 : _GEN_736; // @[CharOutput.scala 82:{21,21}]
  wire [3:0] _GEN_738 = 7'h1e == _char_index_3_T_1[6:0] ? 4'h3 : _GEN_737; // @[CharOutput.scala 82:{21,21}]
  wire [3:0] _GEN_739 = 7'h1f == _char_index_3_T_1[6:0] ? 4'h3 : _GEN_738; // @[CharOutput.scala 82:{21,21}]
  wire [3:0] _GEN_740 = 7'h20 == _char_index_3_T_1[6:0] ? 4'h3 : _GEN_739; // @[CharOutput.scala 82:{21,21}]
  wire [3:0] _GEN_741 = 7'h21 == _char_index_3_T_1[6:0] ? 4'h3 : _GEN_740; // @[CharOutput.scala 82:{21,21}]
  wire [3:0] _GEN_742 = 7'h22 == _char_index_3_T_1[6:0] ? 4'h3 : _GEN_741; // @[CharOutput.scala 82:{21,21}]
  wire [3:0] _GEN_743 = 7'h23 == _char_index_3_T_1[6:0] ? 4'h3 : _GEN_742; // @[CharOutput.scala 82:{21,21}]
  wire [3:0] _GEN_744 = 7'h24 == _char_index_3_T_1[6:0] ? 4'h4 : _GEN_743; // @[CharOutput.scala 82:{21,21}]
  wire [3:0] _GEN_745 = 7'h25 == _char_index_3_T_1[6:0] ? 4'h4 : _GEN_744; // @[CharOutput.scala 82:{21,21}]
  wire [3:0] _GEN_746 = 7'h26 == _char_index_3_T_1[6:0] ? 4'h4 : _GEN_745; // @[CharOutput.scala 82:{21,21}]
  wire [3:0] _GEN_747 = 7'h27 == _char_index_3_T_1[6:0] ? 4'h4 : _GEN_746; // @[CharOutput.scala 82:{21,21}]
  wire [3:0] _GEN_748 = 7'h28 == _char_index_3_T_1[6:0] ? 4'h4 : _GEN_747; // @[CharOutput.scala 82:{21,21}]
  wire [3:0] _GEN_749 = 7'h29 == _char_index_3_T_1[6:0] ? 4'h4 : _GEN_748; // @[CharOutput.scala 82:{21,21}]
  wire [3:0] _GEN_750 = 7'h2a == _char_index_3_T_1[6:0] ? 4'h4 : _GEN_749; // @[CharOutput.scala 82:{21,21}]
  wire [3:0] _GEN_751 = 7'h2b == _char_index_3_T_1[6:0] ? 4'h4 : _GEN_750; // @[CharOutput.scala 82:{21,21}]
  wire [3:0] _GEN_752 = 7'h2c == _char_index_3_T_1[6:0] ? 4'h4 : _GEN_751; // @[CharOutput.scala 82:{21,21}]
  wire [3:0] _GEN_753 = 7'h2d == _char_index_3_T_1[6:0] ? 4'h5 : _GEN_752; // @[CharOutput.scala 82:{21,21}]
  wire [3:0] _GEN_754 = 7'h2e == _char_index_3_T_1[6:0] ? 4'h5 : _GEN_753; // @[CharOutput.scala 82:{21,21}]
  wire [3:0] _GEN_755 = 7'h2f == _char_index_3_T_1[6:0] ? 4'h5 : _GEN_754; // @[CharOutput.scala 82:{21,21}]
  wire [3:0] _GEN_756 = 7'h30 == _char_index_3_T_1[6:0] ? 4'h5 : _GEN_755; // @[CharOutput.scala 82:{21,21}]
  wire [3:0] _GEN_757 = 7'h31 == _char_index_3_T_1[6:0] ? 4'h5 : _GEN_756; // @[CharOutput.scala 82:{21,21}]
  wire [3:0] _GEN_758 = 7'h32 == _char_index_3_T_1[6:0] ? 4'h5 : _GEN_757; // @[CharOutput.scala 82:{21,21}]
  wire [3:0] _GEN_759 = 7'h33 == _char_index_3_T_1[6:0] ? 4'h5 : _GEN_758; // @[CharOutput.scala 82:{21,21}]
  wire [3:0] _GEN_760 = 7'h34 == _char_index_3_T_1[6:0] ? 4'h5 : _GEN_759; // @[CharOutput.scala 82:{21,21}]
  wire [3:0] _GEN_761 = 7'h35 == _char_index_3_T_1[6:0] ? 4'h5 : _GEN_760; // @[CharOutput.scala 82:{21,21}]
  wire [3:0] _GEN_762 = 7'h36 == _char_index_3_T_1[6:0] ? 4'h6 : _GEN_761; // @[CharOutput.scala 82:{21,21}]
  wire [3:0] _GEN_763 = 7'h37 == _char_index_3_T_1[6:0] ? 4'h6 : _GEN_762; // @[CharOutput.scala 82:{21,21}]
  wire [3:0] _GEN_764 = 7'h38 == _char_index_3_T_1[6:0] ? 4'h6 : _GEN_763; // @[CharOutput.scala 82:{21,21}]
  wire [3:0] _GEN_765 = 7'h39 == _char_index_3_T_1[6:0] ? 4'h6 : _GEN_764; // @[CharOutput.scala 82:{21,21}]
  wire [3:0] _GEN_766 = 7'h3a == _char_index_3_T_1[6:0] ? 4'h6 : _GEN_765; // @[CharOutput.scala 82:{21,21}]
  wire [3:0] _GEN_767 = 7'h3b == _char_index_3_T_1[6:0] ? 4'h6 : _GEN_766; // @[CharOutput.scala 82:{21,21}]
  wire [3:0] _GEN_768 = 7'h3c == _char_index_3_T_1[6:0] ? 4'h6 : _GEN_767; // @[CharOutput.scala 82:{21,21}]
  wire [3:0] _GEN_769 = 7'h3d == _char_index_3_T_1[6:0] ? 4'h6 : _GEN_768; // @[CharOutput.scala 82:{21,21}]
  wire [3:0] _GEN_770 = 7'h3e == _char_index_3_T_1[6:0] ? 4'h6 : _GEN_769; // @[CharOutput.scala 82:{21,21}]
  wire [3:0] _GEN_771 = 7'h3f == _char_index_3_T_1[6:0] ? 4'h7 : _GEN_770; // @[CharOutput.scala 82:{21,21}]
  wire [3:0] _GEN_772 = 7'h40 == _char_index_3_T_1[6:0] ? 4'h7 : _GEN_771; // @[CharOutput.scala 82:{21,21}]
  wire [3:0] _GEN_773 = 7'h41 == _char_index_3_T_1[6:0] ? 4'h7 : _GEN_772; // @[CharOutput.scala 82:{21,21}]
  wire [3:0] _GEN_774 = 7'h42 == _char_index_3_T_1[6:0] ? 4'h7 : _GEN_773; // @[CharOutput.scala 82:{21,21}]
  wire [3:0] _GEN_775 = 7'h43 == _char_index_3_T_1[6:0] ? 4'h7 : _GEN_774; // @[CharOutput.scala 82:{21,21}]
  wire [3:0] _GEN_776 = 7'h44 == _char_index_3_T_1[6:0] ? 4'h7 : _GEN_775; // @[CharOutput.scala 82:{21,21}]
  wire [3:0] _GEN_777 = 7'h45 == _char_index_3_T_1[6:0] ? 4'h7 : _GEN_776; // @[CharOutput.scala 82:{21,21}]
  wire [3:0] _GEN_778 = 7'h46 == _char_index_3_T_1[6:0] ? 4'h7 : _GEN_777; // @[CharOutput.scala 82:{21,21}]
  wire [3:0] _GEN_779 = 7'h47 == _char_index_3_T_1[6:0] ? 4'h7 : _GEN_778; // @[CharOutput.scala 82:{21,21}]
  wire [3:0] _GEN_780 = 7'h48 == _char_index_3_T_1[6:0] ? 4'h8 : _GEN_779; // @[CharOutput.scala 82:{21,21}]
  wire [3:0] _GEN_781 = 7'h49 == _char_index_3_T_1[6:0] ? 4'h8 : _GEN_780; // @[CharOutput.scala 82:{21,21}]
  wire [3:0] _GEN_782 = 7'h4a == _char_index_3_T_1[6:0] ? 4'h8 : _GEN_781; // @[CharOutput.scala 82:{21,21}]
  wire [3:0] _GEN_783 = 7'h4b == _char_index_3_T_1[6:0] ? 4'h8 : _GEN_782; // @[CharOutput.scala 82:{21,21}]
  wire [3:0] _GEN_784 = 7'h4c == _char_index_3_T_1[6:0] ? 4'h8 : _GEN_783; // @[CharOutput.scala 82:{21,21}]
  wire [3:0] _GEN_785 = 7'h4d == _char_index_3_T_1[6:0] ? 4'h8 : _GEN_784; // @[CharOutput.scala 82:{21,21}]
  wire [3:0] _GEN_786 = 7'h4e == _char_index_3_T_1[6:0] ? 4'h8 : _GEN_785; // @[CharOutput.scala 82:{21,21}]
  wire [3:0] _GEN_787 = 7'h4f == _char_index_3_T_1[6:0] ? 4'h8 : _GEN_786; // @[CharOutput.scala 82:{21,21}]
  wire [3:0] _GEN_788 = 7'h50 == _char_index_3_T_1[6:0] ? 4'h8 : _GEN_787; // @[CharOutput.scala 82:{21,21}]
  wire [3:0] _GEN_789 = 7'h51 == _char_index_3_T_1[6:0] ? 4'h9 : _GEN_788; // @[CharOutput.scala 82:{21,21}]
  wire [3:0] _GEN_790 = 7'h52 == _char_index_3_T_1[6:0] ? 4'h9 : _GEN_789; // @[CharOutput.scala 82:{21,21}]
  wire [3:0] _GEN_791 = 7'h53 == _char_index_3_T_1[6:0] ? 4'h9 : _GEN_790; // @[CharOutput.scala 82:{21,21}]
  wire [3:0] _GEN_792 = 7'h54 == _char_index_3_T_1[6:0] ? 4'h9 : _GEN_791; // @[CharOutput.scala 82:{21,21}]
  wire [3:0] _GEN_793 = 7'h55 == _char_index_3_T_1[6:0] ? 4'h9 : _GEN_792; // @[CharOutput.scala 82:{21,21}]
  wire [3:0] _GEN_794 = 7'h56 == _char_index_3_T_1[6:0] ? 4'h9 : _GEN_793; // @[CharOutput.scala 82:{21,21}]
  wire [3:0] _GEN_795 = 7'h57 == _char_index_3_T_1[6:0] ? 4'h9 : _GEN_794; // @[CharOutput.scala 82:{21,21}]
  wire [3:0] _GEN_796 = 7'h58 == _char_index_3_T_1[6:0] ? 4'h9 : _GEN_795; // @[CharOutput.scala 82:{21,21}]
  wire [3:0] _GEN_797 = 7'h59 == _char_index_3_T_1[6:0] ? 4'h9 : _GEN_796; // @[CharOutput.scala 82:{21,21}]
  wire [3:0] _GEN_798 = 7'h5a == _char_index_3_T_1[6:0] ? 4'ha : _GEN_797; // @[CharOutput.scala 82:{21,21}]
  wire [3:0] _GEN_799 = 7'h5b == _char_index_3_T_1[6:0] ? 4'ha : _GEN_798; // @[CharOutput.scala 82:{21,21}]
  wire [3:0] _GEN_800 = 7'h5c == _char_index_3_T_1[6:0] ? 4'ha : _GEN_799; // @[CharOutput.scala 82:{21,21}]
  wire [3:0] _GEN_801 = 7'h5d == _char_index_3_T_1[6:0] ? 4'ha : _GEN_800; // @[CharOutput.scala 82:{21,21}]
  wire [3:0] _GEN_802 = 7'h5e == _char_index_3_T_1[6:0] ? 4'ha : _GEN_801; // @[CharOutput.scala 82:{21,21}]
  wire [3:0] _GEN_803 = 7'h5f == _char_index_3_T_1[6:0] ? 4'ha : _GEN_802; // @[CharOutput.scala 82:{21,21}]
  wire [3:0] _GEN_804 = 7'h60 == _char_index_3_T_1[6:0] ? 4'ha : _GEN_803; // @[CharOutput.scala 82:{21,21}]
  wire [3:0] _GEN_805 = 7'h61 == _char_index_3_T_1[6:0] ? 4'ha : _GEN_804; // @[CharOutput.scala 82:{21,21}]
  wire [3:0] _GEN_806 = 7'h62 == _char_index_3_T_1[6:0] ? 4'ha : _GEN_805; // @[CharOutput.scala 82:{21,21}]
  wire [3:0] _GEN_808 = 7'h1 == _char_index_3_T_1[6:0] ? 4'h1 : 4'h0; // @[CharOutput.scala 83:{19,19}]
  wire [3:0] _GEN_809 = 7'h2 == _char_index_3_T_1[6:0] ? 4'h2 : _GEN_808; // @[CharOutput.scala 83:{19,19}]
  wire [3:0] _GEN_810 = 7'h3 == _char_index_3_T_1[6:0] ? 4'h3 : _GEN_809; // @[CharOutput.scala 83:{19,19}]
  wire [3:0] _GEN_811 = 7'h4 == _char_index_3_T_1[6:0] ? 4'h4 : _GEN_810; // @[CharOutput.scala 83:{19,19}]
  wire [3:0] _GEN_812 = 7'h5 == _char_index_3_T_1[6:0] ? 4'h5 : _GEN_811; // @[CharOutput.scala 83:{19,19}]
  wire [3:0] _GEN_813 = 7'h6 == _char_index_3_T_1[6:0] ? 4'h6 : _GEN_812; // @[CharOutput.scala 83:{19,19}]
  wire [3:0] _GEN_814 = 7'h7 == _char_index_3_T_1[6:0] ? 4'h7 : _GEN_813; // @[CharOutput.scala 83:{19,19}]
  wire [3:0] _GEN_815 = 7'h8 == _char_index_3_T_1[6:0] ? 4'h8 : _GEN_814; // @[CharOutput.scala 83:{19,19}]
  wire [3:0] _GEN_816 = 7'h9 == _char_index_3_T_1[6:0] ? 4'h0 : _GEN_815; // @[CharOutput.scala 83:{19,19}]
  wire [3:0] _GEN_817 = 7'ha == _char_index_3_T_1[6:0] ? 4'h1 : _GEN_816; // @[CharOutput.scala 83:{19,19}]
  wire [3:0] _GEN_818 = 7'hb == _char_index_3_T_1[6:0] ? 4'h2 : _GEN_817; // @[CharOutput.scala 83:{19,19}]
  wire [3:0] _GEN_819 = 7'hc == _char_index_3_T_1[6:0] ? 4'h3 : _GEN_818; // @[CharOutput.scala 83:{19,19}]
  wire [3:0] _GEN_820 = 7'hd == _char_index_3_T_1[6:0] ? 4'h4 : _GEN_819; // @[CharOutput.scala 83:{19,19}]
  wire [3:0] _GEN_821 = 7'he == _char_index_3_T_1[6:0] ? 4'h5 : _GEN_820; // @[CharOutput.scala 83:{19,19}]
  wire [3:0] _GEN_822 = 7'hf == _char_index_3_T_1[6:0] ? 4'h6 : _GEN_821; // @[CharOutput.scala 83:{19,19}]
  wire [3:0] _GEN_823 = 7'h10 == _char_index_3_T_1[6:0] ? 4'h7 : _GEN_822; // @[CharOutput.scala 83:{19,19}]
  wire [3:0] _GEN_824 = 7'h11 == _char_index_3_T_1[6:0] ? 4'h8 : _GEN_823; // @[CharOutput.scala 83:{19,19}]
  wire [3:0] _GEN_825 = 7'h12 == _char_index_3_T_1[6:0] ? 4'h0 : _GEN_824; // @[CharOutput.scala 83:{19,19}]
  wire [3:0] _GEN_826 = 7'h13 == _char_index_3_T_1[6:0] ? 4'h1 : _GEN_825; // @[CharOutput.scala 83:{19,19}]
  wire [3:0] _GEN_827 = 7'h14 == _char_index_3_T_1[6:0] ? 4'h2 : _GEN_826; // @[CharOutput.scala 83:{19,19}]
  wire [3:0] _GEN_828 = 7'h15 == _char_index_3_T_1[6:0] ? 4'h3 : _GEN_827; // @[CharOutput.scala 83:{19,19}]
  wire [3:0] _GEN_829 = 7'h16 == _char_index_3_T_1[6:0] ? 4'h4 : _GEN_828; // @[CharOutput.scala 83:{19,19}]
  wire [3:0] _GEN_830 = 7'h17 == _char_index_3_T_1[6:0] ? 4'h5 : _GEN_829; // @[CharOutput.scala 83:{19,19}]
  wire [3:0] _GEN_831 = 7'h18 == _char_index_3_T_1[6:0] ? 4'h6 : _GEN_830; // @[CharOutput.scala 83:{19,19}]
  wire [3:0] _GEN_832 = 7'h19 == _char_index_3_T_1[6:0] ? 4'h7 : _GEN_831; // @[CharOutput.scala 83:{19,19}]
  wire [3:0] _GEN_833 = 7'h1a == _char_index_3_T_1[6:0] ? 4'h8 : _GEN_832; // @[CharOutput.scala 83:{19,19}]
  wire [3:0] _GEN_834 = 7'h1b == _char_index_3_T_1[6:0] ? 4'h0 : _GEN_833; // @[CharOutput.scala 83:{19,19}]
  wire [3:0] _GEN_835 = 7'h1c == _char_index_3_T_1[6:0] ? 4'h1 : _GEN_834; // @[CharOutput.scala 83:{19,19}]
  wire [3:0] _GEN_836 = 7'h1d == _char_index_3_T_1[6:0] ? 4'h2 : _GEN_835; // @[CharOutput.scala 83:{19,19}]
  wire [3:0] _GEN_837 = 7'h1e == _char_index_3_T_1[6:0] ? 4'h3 : _GEN_836; // @[CharOutput.scala 83:{19,19}]
  wire [3:0] _GEN_838 = 7'h1f == _char_index_3_T_1[6:0] ? 4'h4 : _GEN_837; // @[CharOutput.scala 83:{19,19}]
  wire [3:0] _GEN_839 = 7'h20 == _char_index_3_T_1[6:0] ? 4'h5 : _GEN_838; // @[CharOutput.scala 83:{19,19}]
  wire [3:0] _GEN_840 = 7'h21 == _char_index_3_T_1[6:0] ? 4'h6 : _GEN_839; // @[CharOutput.scala 83:{19,19}]
  wire [3:0] _GEN_841 = 7'h22 == _char_index_3_T_1[6:0] ? 4'h7 : _GEN_840; // @[CharOutput.scala 83:{19,19}]
  wire [3:0] _GEN_842 = 7'h23 == _char_index_3_T_1[6:0] ? 4'h8 : _GEN_841; // @[CharOutput.scala 83:{19,19}]
  wire [3:0] _GEN_843 = 7'h24 == _char_index_3_T_1[6:0] ? 4'h0 : _GEN_842; // @[CharOutput.scala 83:{19,19}]
  wire [3:0] _GEN_844 = 7'h25 == _char_index_3_T_1[6:0] ? 4'h1 : _GEN_843; // @[CharOutput.scala 83:{19,19}]
  wire [3:0] _GEN_845 = 7'h26 == _char_index_3_T_1[6:0] ? 4'h2 : _GEN_844; // @[CharOutput.scala 83:{19,19}]
  wire [3:0] _GEN_846 = 7'h27 == _char_index_3_T_1[6:0] ? 4'h3 : _GEN_845; // @[CharOutput.scala 83:{19,19}]
  wire [3:0] _GEN_847 = 7'h28 == _char_index_3_T_1[6:0] ? 4'h4 : _GEN_846; // @[CharOutput.scala 83:{19,19}]
  wire [3:0] _GEN_848 = 7'h29 == _char_index_3_T_1[6:0] ? 4'h5 : _GEN_847; // @[CharOutput.scala 83:{19,19}]
  wire [3:0] _GEN_849 = 7'h2a == _char_index_3_T_1[6:0] ? 4'h6 : _GEN_848; // @[CharOutput.scala 83:{19,19}]
  wire [3:0] _GEN_850 = 7'h2b == _char_index_3_T_1[6:0] ? 4'h7 : _GEN_849; // @[CharOutput.scala 83:{19,19}]
  wire [3:0] _GEN_851 = 7'h2c == _char_index_3_T_1[6:0] ? 4'h8 : _GEN_850; // @[CharOutput.scala 83:{19,19}]
  wire [3:0] _GEN_852 = 7'h2d == _char_index_3_T_1[6:0] ? 4'h0 : _GEN_851; // @[CharOutput.scala 83:{19,19}]
  wire [3:0] _GEN_853 = 7'h2e == _char_index_3_T_1[6:0] ? 4'h1 : _GEN_852; // @[CharOutput.scala 83:{19,19}]
  wire [3:0] _GEN_854 = 7'h2f == _char_index_3_T_1[6:0] ? 4'h2 : _GEN_853; // @[CharOutput.scala 83:{19,19}]
  wire [3:0] _GEN_855 = 7'h30 == _char_index_3_T_1[6:0] ? 4'h3 : _GEN_854; // @[CharOutput.scala 83:{19,19}]
  wire [3:0] _GEN_856 = 7'h31 == _char_index_3_T_1[6:0] ? 4'h4 : _GEN_855; // @[CharOutput.scala 83:{19,19}]
  wire [3:0] _GEN_857 = 7'h32 == _char_index_3_T_1[6:0] ? 4'h5 : _GEN_856; // @[CharOutput.scala 83:{19,19}]
  wire [3:0] _GEN_858 = 7'h33 == _char_index_3_T_1[6:0] ? 4'h6 : _GEN_857; // @[CharOutput.scala 83:{19,19}]
  wire [3:0] _GEN_859 = 7'h34 == _char_index_3_T_1[6:0] ? 4'h7 : _GEN_858; // @[CharOutput.scala 83:{19,19}]
  wire [3:0] _GEN_860 = 7'h35 == _char_index_3_T_1[6:0] ? 4'h8 : _GEN_859; // @[CharOutput.scala 83:{19,19}]
  wire [3:0] _GEN_861 = 7'h36 == _char_index_3_T_1[6:0] ? 4'h0 : _GEN_860; // @[CharOutput.scala 83:{19,19}]
  wire [3:0] _GEN_862 = 7'h37 == _char_index_3_T_1[6:0] ? 4'h1 : _GEN_861; // @[CharOutput.scala 83:{19,19}]
  wire [3:0] _GEN_863 = 7'h38 == _char_index_3_T_1[6:0] ? 4'h2 : _GEN_862; // @[CharOutput.scala 83:{19,19}]
  wire [3:0] _GEN_864 = 7'h39 == _char_index_3_T_1[6:0] ? 4'h3 : _GEN_863; // @[CharOutput.scala 83:{19,19}]
  wire [3:0] _GEN_865 = 7'h3a == _char_index_3_T_1[6:0] ? 4'h4 : _GEN_864; // @[CharOutput.scala 83:{19,19}]
  wire [3:0] _GEN_866 = 7'h3b == _char_index_3_T_1[6:0] ? 4'h5 : _GEN_865; // @[CharOutput.scala 83:{19,19}]
  wire [3:0] _GEN_867 = 7'h3c == _char_index_3_T_1[6:0] ? 4'h6 : _GEN_866; // @[CharOutput.scala 83:{19,19}]
  wire [3:0] _GEN_868 = 7'h3d == _char_index_3_T_1[6:0] ? 4'h7 : _GEN_867; // @[CharOutput.scala 83:{19,19}]
  wire [3:0] _GEN_869 = 7'h3e == _char_index_3_T_1[6:0] ? 4'h8 : _GEN_868; // @[CharOutput.scala 83:{19,19}]
  wire [3:0] _GEN_870 = 7'h3f == _char_index_3_T_1[6:0] ? 4'h0 : _GEN_869; // @[CharOutput.scala 83:{19,19}]
  wire [3:0] _GEN_871 = 7'h40 == _char_index_3_T_1[6:0] ? 4'h1 : _GEN_870; // @[CharOutput.scala 83:{19,19}]
  wire [3:0] _GEN_872 = 7'h41 == _char_index_3_T_1[6:0] ? 4'h2 : _GEN_871; // @[CharOutput.scala 83:{19,19}]
  wire [3:0] _GEN_873 = 7'h42 == _char_index_3_T_1[6:0] ? 4'h3 : _GEN_872; // @[CharOutput.scala 83:{19,19}]
  wire [3:0] _GEN_874 = 7'h43 == _char_index_3_T_1[6:0] ? 4'h4 : _GEN_873; // @[CharOutput.scala 83:{19,19}]
  wire [3:0] _GEN_875 = 7'h44 == _char_index_3_T_1[6:0] ? 4'h5 : _GEN_874; // @[CharOutput.scala 83:{19,19}]
  wire [3:0] _GEN_876 = 7'h45 == _char_index_3_T_1[6:0] ? 4'h6 : _GEN_875; // @[CharOutput.scala 83:{19,19}]
  wire [3:0] _GEN_877 = 7'h46 == _char_index_3_T_1[6:0] ? 4'h7 : _GEN_876; // @[CharOutput.scala 83:{19,19}]
  wire [3:0] _GEN_878 = 7'h47 == _char_index_3_T_1[6:0] ? 4'h8 : _GEN_877; // @[CharOutput.scala 83:{19,19}]
  wire [3:0] _GEN_879 = 7'h48 == _char_index_3_T_1[6:0] ? 4'h0 : _GEN_878; // @[CharOutput.scala 83:{19,19}]
  wire [3:0] _GEN_880 = 7'h49 == _char_index_3_T_1[6:0] ? 4'h1 : _GEN_879; // @[CharOutput.scala 83:{19,19}]
  wire [3:0] _GEN_881 = 7'h4a == _char_index_3_T_1[6:0] ? 4'h2 : _GEN_880; // @[CharOutput.scala 83:{19,19}]
  wire [3:0] _GEN_882 = 7'h4b == _char_index_3_T_1[6:0] ? 4'h3 : _GEN_881; // @[CharOutput.scala 83:{19,19}]
  wire [3:0] _GEN_883 = 7'h4c == _char_index_3_T_1[6:0] ? 4'h4 : _GEN_882; // @[CharOutput.scala 83:{19,19}]
  wire [3:0] _GEN_884 = 7'h4d == _char_index_3_T_1[6:0] ? 4'h5 : _GEN_883; // @[CharOutput.scala 83:{19,19}]
  wire [3:0] _GEN_885 = 7'h4e == _char_index_3_T_1[6:0] ? 4'h6 : _GEN_884; // @[CharOutput.scala 83:{19,19}]
  wire [3:0] _GEN_886 = 7'h4f == _char_index_3_T_1[6:0] ? 4'h7 : _GEN_885; // @[CharOutput.scala 83:{19,19}]
  wire [3:0] _GEN_887 = 7'h50 == _char_index_3_T_1[6:0] ? 4'h8 : _GEN_886; // @[CharOutput.scala 83:{19,19}]
  wire [3:0] _GEN_888 = 7'h51 == _char_index_3_T_1[6:0] ? 4'h0 : _GEN_887; // @[CharOutput.scala 83:{19,19}]
  wire [3:0] _GEN_889 = 7'h52 == _char_index_3_T_1[6:0] ? 4'h1 : _GEN_888; // @[CharOutput.scala 83:{19,19}]
  wire [3:0] _GEN_890 = 7'h53 == _char_index_3_T_1[6:0] ? 4'h2 : _GEN_889; // @[CharOutput.scala 83:{19,19}]
  wire [3:0] _GEN_891 = 7'h54 == _char_index_3_T_1[6:0] ? 4'h3 : _GEN_890; // @[CharOutput.scala 83:{19,19}]
  wire [3:0] _GEN_892 = 7'h55 == _char_index_3_T_1[6:0] ? 4'h4 : _GEN_891; // @[CharOutput.scala 83:{19,19}]
  wire [3:0] _GEN_893 = 7'h56 == _char_index_3_T_1[6:0] ? 4'h5 : _GEN_892; // @[CharOutput.scala 83:{19,19}]
  wire [3:0] _GEN_894 = 7'h57 == _char_index_3_T_1[6:0] ? 4'h6 : _GEN_893; // @[CharOutput.scala 83:{19,19}]
  wire [3:0] _GEN_895 = 7'h58 == _char_index_3_T_1[6:0] ? 4'h7 : _GEN_894; // @[CharOutput.scala 83:{19,19}]
  wire [3:0] _GEN_896 = 7'h59 == _char_index_3_T_1[6:0] ? 4'h8 : _GEN_895; // @[CharOutput.scala 83:{19,19}]
  wire [3:0] _GEN_897 = 7'h5a == _char_index_3_T_1[6:0] ? 4'h0 : _GEN_896; // @[CharOutput.scala 83:{19,19}]
  wire [3:0] _GEN_898 = 7'h5b == _char_index_3_T_1[6:0] ? 4'h1 : _GEN_897; // @[CharOutput.scala 83:{19,19}]
  wire [3:0] _GEN_899 = 7'h5c == _char_index_3_T_1[6:0] ? 4'h2 : _GEN_898; // @[CharOutput.scala 83:{19,19}]
  wire [3:0] _GEN_900 = 7'h5d == _char_index_3_T_1[6:0] ? 4'h3 : _GEN_899; // @[CharOutput.scala 83:{19,19}]
  wire [3:0] _GEN_901 = 7'h5e == _char_index_3_T_1[6:0] ? 4'h4 : _GEN_900; // @[CharOutput.scala 83:{19,19}]
  wire [3:0] _GEN_902 = 7'h5f == _char_index_3_T_1[6:0] ? 4'h5 : _GEN_901; // @[CharOutput.scala 83:{19,19}]
  wire [3:0] _GEN_903 = 7'h60 == _char_index_3_T_1[6:0] ? 4'h6 : _GEN_902; // @[CharOutput.scala 83:{19,19}]
  wire [3:0] _GEN_904 = 7'h61 == _char_index_3_T_1[6:0] ? 4'h7 : _GEN_903; // @[CharOutput.scala 83:{19,19}]
  wire [3:0] _GEN_905 = 7'h62 == _char_index_3_T_1[6:0] ? 4'h8 : _GEN_904; // @[CharOutput.scala 83:{19,19}]
  wire [3:0] char_index_3 = in_area_h_3 ? _GEN_806 : 4'h0; // @[CharOutput.scala 81:23 82:21 85:21]
  wire [3:0] char_col_3 = in_area_h_3 ? _GEN_905 : 4'h0; // @[CharOutput.scala 81:23 83:19 86:19]
  wire [10:0] _char_row_3_T_1 = io_v_cnt - char_area_ytop_3; // @[CharOutput.scala 89:31]
  wire [10:0] _GEN_908 = in_area_v_3 ? _char_row_3_T_1 : 11'h0; // @[CharOutput.scala 88:23 89:19 91:19]
  wire [10:0] _char_index_4_T_1 = io_h_cnt - io_rect_xleft_4; // @[CharOutput.scala 82:48]
  wire [3:0] _GEN_918 = 7'h9 == _char_index_4_T_1[6:0] ? 4'h1 : 4'h0; // @[CharOutput.scala 82:{21,21}]
  wire [3:0] _GEN_919 = 7'ha == _char_index_4_T_1[6:0] ? 4'h1 : _GEN_918; // @[CharOutput.scala 82:{21,21}]
  wire [3:0] _GEN_920 = 7'hb == _char_index_4_T_1[6:0] ? 4'h1 : _GEN_919; // @[CharOutput.scala 82:{21,21}]
  wire [3:0] _GEN_921 = 7'hc == _char_index_4_T_1[6:0] ? 4'h1 : _GEN_920; // @[CharOutput.scala 82:{21,21}]
  wire [3:0] _GEN_922 = 7'hd == _char_index_4_T_1[6:0] ? 4'h1 : _GEN_921; // @[CharOutput.scala 82:{21,21}]
  wire [3:0] _GEN_923 = 7'he == _char_index_4_T_1[6:0] ? 4'h1 : _GEN_922; // @[CharOutput.scala 82:{21,21}]
  wire [3:0] _GEN_924 = 7'hf == _char_index_4_T_1[6:0] ? 4'h1 : _GEN_923; // @[CharOutput.scala 82:{21,21}]
  wire [3:0] _GEN_925 = 7'h10 == _char_index_4_T_1[6:0] ? 4'h1 : _GEN_924; // @[CharOutput.scala 82:{21,21}]
  wire [3:0] _GEN_926 = 7'h11 == _char_index_4_T_1[6:0] ? 4'h1 : _GEN_925; // @[CharOutput.scala 82:{21,21}]
  wire [3:0] _GEN_927 = 7'h12 == _char_index_4_T_1[6:0] ? 4'h2 : _GEN_926; // @[CharOutput.scala 82:{21,21}]
  wire [3:0] _GEN_928 = 7'h13 == _char_index_4_T_1[6:0] ? 4'h2 : _GEN_927; // @[CharOutput.scala 82:{21,21}]
  wire [3:0] _GEN_929 = 7'h14 == _char_index_4_T_1[6:0] ? 4'h2 : _GEN_928; // @[CharOutput.scala 82:{21,21}]
  wire [3:0] _GEN_930 = 7'h15 == _char_index_4_T_1[6:0] ? 4'h2 : _GEN_929; // @[CharOutput.scala 82:{21,21}]
  wire [3:0] _GEN_931 = 7'h16 == _char_index_4_T_1[6:0] ? 4'h2 : _GEN_930; // @[CharOutput.scala 82:{21,21}]
  wire [3:0] _GEN_932 = 7'h17 == _char_index_4_T_1[6:0] ? 4'h2 : _GEN_931; // @[CharOutput.scala 82:{21,21}]
  wire [3:0] _GEN_933 = 7'h18 == _char_index_4_T_1[6:0] ? 4'h2 : _GEN_932; // @[CharOutput.scala 82:{21,21}]
  wire [3:0] _GEN_934 = 7'h19 == _char_index_4_T_1[6:0] ? 4'h2 : _GEN_933; // @[CharOutput.scala 82:{21,21}]
  wire [3:0] _GEN_935 = 7'h1a == _char_index_4_T_1[6:0] ? 4'h2 : _GEN_934; // @[CharOutput.scala 82:{21,21}]
  wire [3:0] _GEN_936 = 7'h1b == _char_index_4_T_1[6:0] ? 4'h3 : _GEN_935; // @[CharOutput.scala 82:{21,21}]
  wire [3:0] _GEN_937 = 7'h1c == _char_index_4_T_1[6:0] ? 4'h3 : _GEN_936; // @[CharOutput.scala 82:{21,21}]
  wire [3:0] _GEN_938 = 7'h1d == _char_index_4_T_1[6:0] ? 4'h3 : _GEN_937; // @[CharOutput.scala 82:{21,21}]
  wire [3:0] _GEN_939 = 7'h1e == _char_index_4_T_1[6:0] ? 4'h3 : _GEN_938; // @[CharOutput.scala 82:{21,21}]
  wire [3:0] _GEN_940 = 7'h1f == _char_index_4_T_1[6:0] ? 4'h3 : _GEN_939; // @[CharOutput.scala 82:{21,21}]
  wire [3:0] _GEN_941 = 7'h20 == _char_index_4_T_1[6:0] ? 4'h3 : _GEN_940; // @[CharOutput.scala 82:{21,21}]
  wire [3:0] _GEN_942 = 7'h21 == _char_index_4_T_1[6:0] ? 4'h3 : _GEN_941; // @[CharOutput.scala 82:{21,21}]
  wire [3:0] _GEN_943 = 7'h22 == _char_index_4_T_1[6:0] ? 4'h3 : _GEN_942; // @[CharOutput.scala 82:{21,21}]
  wire [3:0] _GEN_944 = 7'h23 == _char_index_4_T_1[6:0] ? 4'h3 : _GEN_943; // @[CharOutput.scala 82:{21,21}]
  wire [3:0] _GEN_945 = 7'h24 == _char_index_4_T_1[6:0] ? 4'h4 : _GEN_944; // @[CharOutput.scala 82:{21,21}]
  wire [3:0] _GEN_946 = 7'h25 == _char_index_4_T_1[6:0] ? 4'h4 : _GEN_945; // @[CharOutput.scala 82:{21,21}]
  wire [3:0] _GEN_947 = 7'h26 == _char_index_4_T_1[6:0] ? 4'h4 : _GEN_946; // @[CharOutput.scala 82:{21,21}]
  wire [3:0] _GEN_948 = 7'h27 == _char_index_4_T_1[6:0] ? 4'h4 : _GEN_947; // @[CharOutput.scala 82:{21,21}]
  wire [3:0] _GEN_949 = 7'h28 == _char_index_4_T_1[6:0] ? 4'h4 : _GEN_948; // @[CharOutput.scala 82:{21,21}]
  wire [3:0] _GEN_950 = 7'h29 == _char_index_4_T_1[6:0] ? 4'h4 : _GEN_949; // @[CharOutput.scala 82:{21,21}]
  wire [3:0] _GEN_951 = 7'h2a == _char_index_4_T_1[6:0] ? 4'h4 : _GEN_950; // @[CharOutput.scala 82:{21,21}]
  wire [3:0] _GEN_952 = 7'h2b == _char_index_4_T_1[6:0] ? 4'h4 : _GEN_951; // @[CharOutput.scala 82:{21,21}]
  wire [3:0] _GEN_953 = 7'h2c == _char_index_4_T_1[6:0] ? 4'h4 : _GEN_952; // @[CharOutput.scala 82:{21,21}]
  wire [3:0] _GEN_954 = 7'h2d == _char_index_4_T_1[6:0] ? 4'h5 : _GEN_953; // @[CharOutput.scala 82:{21,21}]
  wire [3:0] _GEN_955 = 7'h2e == _char_index_4_T_1[6:0] ? 4'h5 : _GEN_954; // @[CharOutput.scala 82:{21,21}]
  wire [3:0] _GEN_956 = 7'h2f == _char_index_4_T_1[6:0] ? 4'h5 : _GEN_955; // @[CharOutput.scala 82:{21,21}]
  wire [3:0] _GEN_957 = 7'h30 == _char_index_4_T_1[6:0] ? 4'h5 : _GEN_956; // @[CharOutput.scala 82:{21,21}]
  wire [3:0] _GEN_958 = 7'h31 == _char_index_4_T_1[6:0] ? 4'h5 : _GEN_957; // @[CharOutput.scala 82:{21,21}]
  wire [3:0] _GEN_959 = 7'h32 == _char_index_4_T_1[6:0] ? 4'h5 : _GEN_958; // @[CharOutput.scala 82:{21,21}]
  wire [3:0] _GEN_960 = 7'h33 == _char_index_4_T_1[6:0] ? 4'h5 : _GEN_959; // @[CharOutput.scala 82:{21,21}]
  wire [3:0] _GEN_961 = 7'h34 == _char_index_4_T_1[6:0] ? 4'h5 : _GEN_960; // @[CharOutput.scala 82:{21,21}]
  wire [3:0] _GEN_962 = 7'h35 == _char_index_4_T_1[6:0] ? 4'h5 : _GEN_961; // @[CharOutput.scala 82:{21,21}]
  wire [3:0] _GEN_963 = 7'h36 == _char_index_4_T_1[6:0] ? 4'h6 : _GEN_962; // @[CharOutput.scala 82:{21,21}]
  wire [3:0] _GEN_964 = 7'h37 == _char_index_4_T_1[6:0] ? 4'h6 : _GEN_963; // @[CharOutput.scala 82:{21,21}]
  wire [3:0] _GEN_965 = 7'h38 == _char_index_4_T_1[6:0] ? 4'h6 : _GEN_964; // @[CharOutput.scala 82:{21,21}]
  wire [3:0] _GEN_966 = 7'h39 == _char_index_4_T_1[6:0] ? 4'h6 : _GEN_965; // @[CharOutput.scala 82:{21,21}]
  wire [3:0] _GEN_967 = 7'h3a == _char_index_4_T_1[6:0] ? 4'h6 : _GEN_966; // @[CharOutput.scala 82:{21,21}]
  wire [3:0] _GEN_968 = 7'h3b == _char_index_4_T_1[6:0] ? 4'h6 : _GEN_967; // @[CharOutput.scala 82:{21,21}]
  wire [3:0] _GEN_969 = 7'h3c == _char_index_4_T_1[6:0] ? 4'h6 : _GEN_968; // @[CharOutput.scala 82:{21,21}]
  wire [3:0] _GEN_970 = 7'h3d == _char_index_4_T_1[6:0] ? 4'h6 : _GEN_969; // @[CharOutput.scala 82:{21,21}]
  wire [3:0] _GEN_971 = 7'h3e == _char_index_4_T_1[6:0] ? 4'h6 : _GEN_970; // @[CharOutput.scala 82:{21,21}]
  wire [3:0] _GEN_972 = 7'h3f == _char_index_4_T_1[6:0] ? 4'h7 : _GEN_971; // @[CharOutput.scala 82:{21,21}]
  wire [3:0] _GEN_973 = 7'h40 == _char_index_4_T_1[6:0] ? 4'h7 : _GEN_972; // @[CharOutput.scala 82:{21,21}]
  wire [3:0] _GEN_974 = 7'h41 == _char_index_4_T_1[6:0] ? 4'h7 : _GEN_973; // @[CharOutput.scala 82:{21,21}]
  wire [3:0] _GEN_975 = 7'h42 == _char_index_4_T_1[6:0] ? 4'h7 : _GEN_974; // @[CharOutput.scala 82:{21,21}]
  wire [3:0] _GEN_976 = 7'h43 == _char_index_4_T_1[6:0] ? 4'h7 : _GEN_975; // @[CharOutput.scala 82:{21,21}]
  wire [3:0] _GEN_977 = 7'h44 == _char_index_4_T_1[6:0] ? 4'h7 : _GEN_976; // @[CharOutput.scala 82:{21,21}]
  wire [3:0] _GEN_978 = 7'h45 == _char_index_4_T_1[6:0] ? 4'h7 : _GEN_977; // @[CharOutput.scala 82:{21,21}]
  wire [3:0] _GEN_979 = 7'h46 == _char_index_4_T_1[6:0] ? 4'h7 : _GEN_978; // @[CharOutput.scala 82:{21,21}]
  wire [3:0] _GEN_980 = 7'h47 == _char_index_4_T_1[6:0] ? 4'h7 : _GEN_979; // @[CharOutput.scala 82:{21,21}]
  wire [3:0] _GEN_981 = 7'h48 == _char_index_4_T_1[6:0] ? 4'h8 : _GEN_980; // @[CharOutput.scala 82:{21,21}]
  wire [3:0] _GEN_982 = 7'h49 == _char_index_4_T_1[6:0] ? 4'h8 : _GEN_981; // @[CharOutput.scala 82:{21,21}]
  wire [3:0] _GEN_983 = 7'h4a == _char_index_4_T_1[6:0] ? 4'h8 : _GEN_982; // @[CharOutput.scala 82:{21,21}]
  wire [3:0] _GEN_984 = 7'h4b == _char_index_4_T_1[6:0] ? 4'h8 : _GEN_983; // @[CharOutput.scala 82:{21,21}]
  wire [3:0] _GEN_985 = 7'h4c == _char_index_4_T_1[6:0] ? 4'h8 : _GEN_984; // @[CharOutput.scala 82:{21,21}]
  wire [3:0] _GEN_986 = 7'h4d == _char_index_4_T_1[6:0] ? 4'h8 : _GEN_985; // @[CharOutput.scala 82:{21,21}]
  wire [3:0] _GEN_987 = 7'h4e == _char_index_4_T_1[6:0] ? 4'h8 : _GEN_986; // @[CharOutput.scala 82:{21,21}]
  wire [3:0] _GEN_988 = 7'h4f == _char_index_4_T_1[6:0] ? 4'h8 : _GEN_987; // @[CharOutput.scala 82:{21,21}]
  wire [3:0] _GEN_989 = 7'h50 == _char_index_4_T_1[6:0] ? 4'h8 : _GEN_988; // @[CharOutput.scala 82:{21,21}]
  wire [3:0] _GEN_990 = 7'h51 == _char_index_4_T_1[6:0] ? 4'h9 : _GEN_989; // @[CharOutput.scala 82:{21,21}]
  wire [3:0] _GEN_991 = 7'h52 == _char_index_4_T_1[6:0] ? 4'h9 : _GEN_990; // @[CharOutput.scala 82:{21,21}]
  wire [3:0] _GEN_992 = 7'h53 == _char_index_4_T_1[6:0] ? 4'h9 : _GEN_991; // @[CharOutput.scala 82:{21,21}]
  wire [3:0] _GEN_993 = 7'h54 == _char_index_4_T_1[6:0] ? 4'h9 : _GEN_992; // @[CharOutput.scala 82:{21,21}]
  wire [3:0] _GEN_994 = 7'h55 == _char_index_4_T_1[6:0] ? 4'h9 : _GEN_993; // @[CharOutput.scala 82:{21,21}]
  wire [3:0] _GEN_995 = 7'h56 == _char_index_4_T_1[6:0] ? 4'h9 : _GEN_994; // @[CharOutput.scala 82:{21,21}]
  wire [3:0] _GEN_996 = 7'h57 == _char_index_4_T_1[6:0] ? 4'h9 : _GEN_995; // @[CharOutput.scala 82:{21,21}]
  wire [3:0] _GEN_997 = 7'h58 == _char_index_4_T_1[6:0] ? 4'h9 : _GEN_996; // @[CharOutput.scala 82:{21,21}]
  wire [3:0] _GEN_998 = 7'h59 == _char_index_4_T_1[6:0] ? 4'h9 : _GEN_997; // @[CharOutput.scala 82:{21,21}]
  wire [3:0] _GEN_999 = 7'h5a == _char_index_4_T_1[6:0] ? 4'ha : _GEN_998; // @[CharOutput.scala 82:{21,21}]
  wire [3:0] _GEN_1000 = 7'h5b == _char_index_4_T_1[6:0] ? 4'ha : _GEN_999; // @[CharOutput.scala 82:{21,21}]
  wire [3:0] _GEN_1001 = 7'h5c == _char_index_4_T_1[6:0] ? 4'ha : _GEN_1000; // @[CharOutput.scala 82:{21,21}]
  wire [3:0] _GEN_1002 = 7'h5d == _char_index_4_T_1[6:0] ? 4'ha : _GEN_1001; // @[CharOutput.scala 82:{21,21}]
  wire [3:0] _GEN_1003 = 7'h5e == _char_index_4_T_1[6:0] ? 4'ha : _GEN_1002; // @[CharOutput.scala 82:{21,21}]
  wire [3:0] _GEN_1004 = 7'h5f == _char_index_4_T_1[6:0] ? 4'ha : _GEN_1003; // @[CharOutput.scala 82:{21,21}]
  wire [3:0] _GEN_1005 = 7'h60 == _char_index_4_T_1[6:0] ? 4'ha : _GEN_1004; // @[CharOutput.scala 82:{21,21}]
  wire [3:0] _GEN_1006 = 7'h61 == _char_index_4_T_1[6:0] ? 4'ha : _GEN_1005; // @[CharOutput.scala 82:{21,21}]
  wire [3:0] _GEN_1007 = 7'h62 == _char_index_4_T_1[6:0] ? 4'ha : _GEN_1006; // @[CharOutput.scala 82:{21,21}]
  wire [3:0] _GEN_1009 = 7'h1 == _char_index_4_T_1[6:0] ? 4'h1 : 4'h0; // @[CharOutput.scala 83:{19,19}]
  wire [3:0] _GEN_1010 = 7'h2 == _char_index_4_T_1[6:0] ? 4'h2 : _GEN_1009; // @[CharOutput.scala 83:{19,19}]
  wire [3:0] _GEN_1011 = 7'h3 == _char_index_4_T_1[6:0] ? 4'h3 : _GEN_1010; // @[CharOutput.scala 83:{19,19}]
  wire [3:0] _GEN_1012 = 7'h4 == _char_index_4_T_1[6:0] ? 4'h4 : _GEN_1011; // @[CharOutput.scala 83:{19,19}]
  wire [3:0] _GEN_1013 = 7'h5 == _char_index_4_T_1[6:0] ? 4'h5 : _GEN_1012; // @[CharOutput.scala 83:{19,19}]
  wire [3:0] _GEN_1014 = 7'h6 == _char_index_4_T_1[6:0] ? 4'h6 : _GEN_1013; // @[CharOutput.scala 83:{19,19}]
  wire [3:0] _GEN_1015 = 7'h7 == _char_index_4_T_1[6:0] ? 4'h7 : _GEN_1014; // @[CharOutput.scala 83:{19,19}]
  wire [3:0] _GEN_1016 = 7'h8 == _char_index_4_T_1[6:0] ? 4'h8 : _GEN_1015; // @[CharOutput.scala 83:{19,19}]
  wire [3:0] _GEN_1017 = 7'h9 == _char_index_4_T_1[6:0] ? 4'h0 : _GEN_1016; // @[CharOutput.scala 83:{19,19}]
  wire [3:0] _GEN_1018 = 7'ha == _char_index_4_T_1[6:0] ? 4'h1 : _GEN_1017; // @[CharOutput.scala 83:{19,19}]
  wire [3:0] _GEN_1019 = 7'hb == _char_index_4_T_1[6:0] ? 4'h2 : _GEN_1018; // @[CharOutput.scala 83:{19,19}]
  wire [3:0] _GEN_1020 = 7'hc == _char_index_4_T_1[6:0] ? 4'h3 : _GEN_1019; // @[CharOutput.scala 83:{19,19}]
  wire [3:0] _GEN_1021 = 7'hd == _char_index_4_T_1[6:0] ? 4'h4 : _GEN_1020; // @[CharOutput.scala 83:{19,19}]
  wire [3:0] _GEN_1022 = 7'he == _char_index_4_T_1[6:0] ? 4'h5 : _GEN_1021; // @[CharOutput.scala 83:{19,19}]
  wire [3:0] _GEN_1023 = 7'hf == _char_index_4_T_1[6:0] ? 4'h6 : _GEN_1022; // @[CharOutput.scala 83:{19,19}]
  wire [3:0] _GEN_1024 = 7'h10 == _char_index_4_T_1[6:0] ? 4'h7 : _GEN_1023; // @[CharOutput.scala 83:{19,19}]
  wire [3:0] _GEN_1025 = 7'h11 == _char_index_4_T_1[6:0] ? 4'h8 : _GEN_1024; // @[CharOutput.scala 83:{19,19}]
  wire [3:0] _GEN_1026 = 7'h12 == _char_index_4_T_1[6:0] ? 4'h0 : _GEN_1025; // @[CharOutput.scala 83:{19,19}]
  wire [3:0] _GEN_1027 = 7'h13 == _char_index_4_T_1[6:0] ? 4'h1 : _GEN_1026; // @[CharOutput.scala 83:{19,19}]
  wire [3:0] _GEN_1028 = 7'h14 == _char_index_4_T_1[6:0] ? 4'h2 : _GEN_1027; // @[CharOutput.scala 83:{19,19}]
  wire [3:0] _GEN_1029 = 7'h15 == _char_index_4_T_1[6:0] ? 4'h3 : _GEN_1028; // @[CharOutput.scala 83:{19,19}]
  wire [3:0] _GEN_1030 = 7'h16 == _char_index_4_T_1[6:0] ? 4'h4 : _GEN_1029; // @[CharOutput.scala 83:{19,19}]
  wire [3:0] _GEN_1031 = 7'h17 == _char_index_4_T_1[6:0] ? 4'h5 : _GEN_1030; // @[CharOutput.scala 83:{19,19}]
  wire [3:0] _GEN_1032 = 7'h18 == _char_index_4_T_1[6:0] ? 4'h6 : _GEN_1031; // @[CharOutput.scala 83:{19,19}]
  wire [3:0] _GEN_1033 = 7'h19 == _char_index_4_T_1[6:0] ? 4'h7 : _GEN_1032; // @[CharOutput.scala 83:{19,19}]
  wire [3:0] _GEN_1034 = 7'h1a == _char_index_4_T_1[6:0] ? 4'h8 : _GEN_1033; // @[CharOutput.scala 83:{19,19}]
  wire [3:0] _GEN_1035 = 7'h1b == _char_index_4_T_1[6:0] ? 4'h0 : _GEN_1034; // @[CharOutput.scala 83:{19,19}]
  wire [3:0] _GEN_1036 = 7'h1c == _char_index_4_T_1[6:0] ? 4'h1 : _GEN_1035; // @[CharOutput.scala 83:{19,19}]
  wire [3:0] _GEN_1037 = 7'h1d == _char_index_4_T_1[6:0] ? 4'h2 : _GEN_1036; // @[CharOutput.scala 83:{19,19}]
  wire [3:0] _GEN_1038 = 7'h1e == _char_index_4_T_1[6:0] ? 4'h3 : _GEN_1037; // @[CharOutput.scala 83:{19,19}]
  wire [3:0] _GEN_1039 = 7'h1f == _char_index_4_T_1[6:0] ? 4'h4 : _GEN_1038; // @[CharOutput.scala 83:{19,19}]
  wire [3:0] _GEN_1040 = 7'h20 == _char_index_4_T_1[6:0] ? 4'h5 : _GEN_1039; // @[CharOutput.scala 83:{19,19}]
  wire [3:0] _GEN_1041 = 7'h21 == _char_index_4_T_1[6:0] ? 4'h6 : _GEN_1040; // @[CharOutput.scala 83:{19,19}]
  wire [3:0] _GEN_1042 = 7'h22 == _char_index_4_T_1[6:0] ? 4'h7 : _GEN_1041; // @[CharOutput.scala 83:{19,19}]
  wire [3:0] _GEN_1043 = 7'h23 == _char_index_4_T_1[6:0] ? 4'h8 : _GEN_1042; // @[CharOutput.scala 83:{19,19}]
  wire [3:0] _GEN_1044 = 7'h24 == _char_index_4_T_1[6:0] ? 4'h0 : _GEN_1043; // @[CharOutput.scala 83:{19,19}]
  wire [3:0] _GEN_1045 = 7'h25 == _char_index_4_T_1[6:0] ? 4'h1 : _GEN_1044; // @[CharOutput.scala 83:{19,19}]
  wire [3:0] _GEN_1046 = 7'h26 == _char_index_4_T_1[6:0] ? 4'h2 : _GEN_1045; // @[CharOutput.scala 83:{19,19}]
  wire [3:0] _GEN_1047 = 7'h27 == _char_index_4_T_1[6:0] ? 4'h3 : _GEN_1046; // @[CharOutput.scala 83:{19,19}]
  wire [3:0] _GEN_1048 = 7'h28 == _char_index_4_T_1[6:0] ? 4'h4 : _GEN_1047; // @[CharOutput.scala 83:{19,19}]
  wire [3:0] _GEN_1049 = 7'h29 == _char_index_4_T_1[6:0] ? 4'h5 : _GEN_1048; // @[CharOutput.scala 83:{19,19}]
  wire [3:0] _GEN_1050 = 7'h2a == _char_index_4_T_1[6:0] ? 4'h6 : _GEN_1049; // @[CharOutput.scala 83:{19,19}]
  wire [3:0] _GEN_1051 = 7'h2b == _char_index_4_T_1[6:0] ? 4'h7 : _GEN_1050; // @[CharOutput.scala 83:{19,19}]
  wire [3:0] _GEN_1052 = 7'h2c == _char_index_4_T_1[6:0] ? 4'h8 : _GEN_1051; // @[CharOutput.scala 83:{19,19}]
  wire [3:0] _GEN_1053 = 7'h2d == _char_index_4_T_1[6:0] ? 4'h0 : _GEN_1052; // @[CharOutput.scala 83:{19,19}]
  wire [3:0] _GEN_1054 = 7'h2e == _char_index_4_T_1[6:0] ? 4'h1 : _GEN_1053; // @[CharOutput.scala 83:{19,19}]
  wire [3:0] _GEN_1055 = 7'h2f == _char_index_4_T_1[6:0] ? 4'h2 : _GEN_1054; // @[CharOutput.scala 83:{19,19}]
  wire [3:0] _GEN_1056 = 7'h30 == _char_index_4_T_1[6:0] ? 4'h3 : _GEN_1055; // @[CharOutput.scala 83:{19,19}]
  wire [3:0] _GEN_1057 = 7'h31 == _char_index_4_T_1[6:0] ? 4'h4 : _GEN_1056; // @[CharOutput.scala 83:{19,19}]
  wire [3:0] _GEN_1058 = 7'h32 == _char_index_4_T_1[6:0] ? 4'h5 : _GEN_1057; // @[CharOutput.scala 83:{19,19}]
  wire [3:0] _GEN_1059 = 7'h33 == _char_index_4_T_1[6:0] ? 4'h6 : _GEN_1058; // @[CharOutput.scala 83:{19,19}]
  wire [3:0] _GEN_1060 = 7'h34 == _char_index_4_T_1[6:0] ? 4'h7 : _GEN_1059; // @[CharOutput.scala 83:{19,19}]
  wire [3:0] _GEN_1061 = 7'h35 == _char_index_4_T_1[6:0] ? 4'h8 : _GEN_1060; // @[CharOutput.scala 83:{19,19}]
  wire [3:0] _GEN_1062 = 7'h36 == _char_index_4_T_1[6:0] ? 4'h0 : _GEN_1061; // @[CharOutput.scala 83:{19,19}]
  wire [3:0] _GEN_1063 = 7'h37 == _char_index_4_T_1[6:0] ? 4'h1 : _GEN_1062; // @[CharOutput.scala 83:{19,19}]
  wire [3:0] _GEN_1064 = 7'h38 == _char_index_4_T_1[6:0] ? 4'h2 : _GEN_1063; // @[CharOutput.scala 83:{19,19}]
  wire [3:0] _GEN_1065 = 7'h39 == _char_index_4_T_1[6:0] ? 4'h3 : _GEN_1064; // @[CharOutput.scala 83:{19,19}]
  wire [3:0] _GEN_1066 = 7'h3a == _char_index_4_T_1[6:0] ? 4'h4 : _GEN_1065; // @[CharOutput.scala 83:{19,19}]
  wire [3:0] _GEN_1067 = 7'h3b == _char_index_4_T_1[6:0] ? 4'h5 : _GEN_1066; // @[CharOutput.scala 83:{19,19}]
  wire [3:0] _GEN_1068 = 7'h3c == _char_index_4_T_1[6:0] ? 4'h6 : _GEN_1067; // @[CharOutput.scala 83:{19,19}]
  wire [3:0] _GEN_1069 = 7'h3d == _char_index_4_T_1[6:0] ? 4'h7 : _GEN_1068; // @[CharOutput.scala 83:{19,19}]
  wire [3:0] _GEN_1070 = 7'h3e == _char_index_4_T_1[6:0] ? 4'h8 : _GEN_1069; // @[CharOutput.scala 83:{19,19}]
  wire [3:0] _GEN_1071 = 7'h3f == _char_index_4_T_1[6:0] ? 4'h0 : _GEN_1070; // @[CharOutput.scala 83:{19,19}]
  wire [3:0] _GEN_1072 = 7'h40 == _char_index_4_T_1[6:0] ? 4'h1 : _GEN_1071; // @[CharOutput.scala 83:{19,19}]
  wire [3:0] _GEN_1073 = 7'h41 == _char_index_4_T_1[6:0] ? 4'h2 : _GEN_1072; // @[CharOutput.scala 83:{19,19}]
  wire [3:0] _GEN_1074 = 7'h42 == _char_index_4_T_1[6:0] ? 4'h3 : _GEN_1073; // @[CharOutput.scala 83:{19,19}]
  wire [3:0] _GEN_1075 = 7'h43 == _char_index_4_T_1[6:0] ? 4'h4 : _GEN_1074; // @[CharOutput.scala 83:{19,19}]
  wire [3:0] _GEN_1076 = 7'h44 == _char_index_4_T_1[6:0] ? 4'h5 : _GEN_1075; // @[CharOutput.scala 83:{19,19}]
  wire [3:0] _GEN_1077 = 7'h45 == _char_index_4_T_1[6:0] ? 4'h6 : _GEN_1076; // @[CharOutput.scala 83:{19,19}]
  wire [3:0] _GEN_1078 = 7'h46 == _char_index_4_T_1[6:0] ? 4'h7 : _GEN_1077; // @[CharOutput.scala 83:{19,19}]
  wire [3:0] _GEN_1079 = 7'h47 == _char_index_4_T_1[6:0] ? 4'h8 : _GEN_1078; // @[CharOutput.scala 83:{19,19}]
  wire [3:0] _GEN_1080 = 7'h48 == _char_index_4_T_1[6:0] ? 4'h0 : _GEN_1079; // @[CharOutput.scala 83:{19,19}]
  wire [3:0] _GEN_1081 = 7'h49 == _char_index_4_T_1[6:0] ? 4'h1 : _GEN_1080; // @[CharOutput.scala 83:{19,19}]
  wire [3:0] _GEN_1082 = 7'h4a == _char_index_4_T_1[6:0] ? 4'h2 : _GEN_1081; // @[CharOutput.scala 83:{19,19}]
  wire [3:0] _GEN_1083 = 7'h4b == _char_index_4_T_1[6:0] ? 4'h3 : _GEN_1082; // @[CharOutput.scala 83:{19,19}]
  wire [3:0] _GEN_1084 = 7'h4c == _char_index_4_T_1[6:0] ? 4'h4 : _GEN_1083; // @[CharOutput.scala 83:{19,19}]
  wire [3:0] _GEN_1085 = 7'h4d == _char_index_4_T_1[6:0] ? 4'h5 : _GEN_1084; // @[CharOutput.scala 83:{19,19}]
  wire [3:0] _GEN_1086 = 7'h4e == _char_index_4_T_1[6:0] ? 4'h6 : _GEN_1085; // @[CharOutput.scala 83:{19,19}]
  wire [3:0] _GEN_1087 = 7'h4f == _char_index_4_T_1[6:0] ? 4'h7 : _GEN_1086; // @[CharOutput.scala 83:{19,19}]
  wire [3:0] _GEN_1088 = 7'h50 == _char_index_4_T_1[6:0] ? 4'h8 : _GEN_1087; // @[CharOutput.scala 83:{19,19}]
  wire [3:0] _GEN_1089 = 7'h51 == _char_index_4_T_1[6:0] ? 4'h0 : _GEN_1088; // @[CharOutput.scala 83:{19,19}]
  wire [3:0] _GEN_1090 = 7'h52 == _char_index_4_T_1[6:0] ? 4'h1 : _GEN_1089; // @[CharOutput.scala 83:{19,19}]
  wire [3:0] _GEN_1091 = 7'h53 == _char_index_4_T_1[6:0] ? 4'h2 : _GEN_1090; // @[CharOutput.scala 83:{19,19}]
  wire [3:0] _GEN_1092 = 7'h54 == _char_index_4_T_1[6:0] ? 4'h3 : _GEN_1091; // @[CharOutput.scala 83:{19,19}]
  wire [3:0] _GEN_1093 = 7'h55 == _char_index_4_T_1[6:0] ? 4'h4 : _GEN_1092; // @[CharOutput.scala 83:{19,19}]
  wire [3:0] _GEN_1094 = 7'h56 == _char_index_4_T_1[6:0] ? 4'h5 : _GEN_1093; // @[CharOutput.scala 83:{19,19}]
  wire [3:0] _GEN_1095 = 7'h57 == _char_index_4_T_1[6:0] ? 4'h6 : _GEN_1094; // @[CharOutput.scala 83:{19,19}]
  wire [3:0] _GEN_1096 = 7'h58 == _char_index_4_T_1[6:0] ? 4'h7 : _GEN_1095; // @[CharOutput.scala 83:{19,19}]
  wire [3:0] _GEN_1097 = 7'h59 == _char_index_4_T_1[6:0] ? 4'h8 : _GEN_1096; // @[CharOutput.scala 83:{19,19}]
  wire [3:0] _GEN_1098 = 7'h5a == _char_index_4_T_1[6:0] ? 4'h0 : _GEN_1097; // @[CharOutput.scala 83:{19,19}]
  wire [3:0] _GEN_1099 = 7'h5b == _char_index_4_T_1[6:0] ? 4'h1 : _GEN_1098; // @[CharOutput.scala 83:{19,19}]
  wire [3:0] _GEN_1100 = 7'h5c == _char_index_4_T_1[6:0] ? 4'h2 : _GEN_1099; // @[CharOutput.scala 83:{19,19}]
  wire [3:0] _GEN_1101 = 7'h5d == _char_index_4_T_1[6:0] ? 4'h3 : _GEN_1100; // @[CharOutput.scala 83:{19,19}]
  wire [3:0] _GEN_1102 = 7'h5e == _char_index_4_T_1[6:0] ? 4'h4 : _GEN_1101; // @[CharOutput.scala 83:{19,19}]
  wire [3:0] _GEN_1103 = 7'h5f == _char_index_4_T_1[6:0] ? 4'h5 : _GEN_1102; // @[CharOutput.scala 83:{19,19}]
  wire [3:0] _GEN_1104 = 7'h60 == _char_index_4_T_1[6:0] ? 4'h6 : _GEN_1103; // @[CharOutput.scala 83:{19,19}]
  wire [3:0] _GEN_1105 = 7'h61 == _char_index_4_T_1[6:0] ? 4'h7 : _GEN_1104; // @[CharOutput.scala 83:{19,19}]
  wire [3:0] _GEN_1106 = 7'h62 == _char_index_4_T_1[6:0] ? 4'h8 : _GEN_1105; // @[CharOutput.scala 83:{19,19}]
  wire [3:0] char_index_4 = in_area_h_4 ? _GEN_1007 : 4'h0; // @[CharOutput.scala 81:23 82:21 85:21]
  wire [3:0] char_col_4 = in_area_h_4 ? _GEN_1106 : 4'h0; // @[CharOutput.scala 81:23 83:19 86:19]
  wire [10:0] _char_row_4_T_1 = io_v_cnt - char_area_ytop_4; // @[CharOutput.scala 89:31]
  wire [10:0] _GEN_1109 = in_area_v_4 ? _char_row_4_T_1 : 11'h0; // @[CharOutput.scala 88:23 89:19 91:19]
  wire  _T_11 = ~char_area_valid_5; // @[CharOutput.scala 98:8]
  wire [2:0] _obj_choose_T = char_area_en_4 ? 3'h4 : 3'h5; // @[Mux.scala 47:70]
  wire [2:0] _obj_choose_T_1 = char_area_en_3 ? 3'h3 : _obj_choose_T; // @[Mux.scala 47:70]
  wire [2:0] _obj_choose_T_2 = char_area_en_2 ? 3'h2 : _obj_choose_T_1; // @[Mux.scala 47:70]
  wire [2:0] _obj_choose_T_3 = char_area_en_1 ? 3'h1 : _obj_choose_T_2; // @[Mux.scala 47:70]
  wire [2:0] _obj_choose_T_4 = char_area_en_0 ? 3'h0 : _obj_choose_T_3; // @[Mux.scala 47:70]
  wire [2:0] obj_choose = ~char_area_valid_5 ? _obj_choose_T_4 : 3'h0; // @[CharOutput.scala 101:16 98:34 99:16]
  wire [5:0] _char_baseaddr_lut_T = 1'h0 * 5'h10; // @[CharOutput.scala 110:60]
  wire [5:0] _char_baseaddr_lut_T_1 = 1'h1 * 5'h10; // @[CharOutput.scala 110:60]
  wire [6:0] _char_baseaddr_lut_T_2 = 2'h2 * 5'h10; // @[CharOutput.scala 110:60]
  wire [6:0] _char_baseaddr_lut_T_3 = 2'h3 * 5'h10; // @[CharOutput.scala 110:60]
  wire [7:0] _char_baseaddr_lut_T_4 = 3'h4 * 5'h10; // @[CharOutput.scala 110:60]
  wire [7:0] _char_baseaddr_lut_T_5 = 3'h5 * 5'h10; // @[CharOutput.scala 110:60]
  wire [7:0] _char_baseaddr_lut_T_6 = 3'h6 * 5'h10; // @[CharOutput.scala 110:60]
  wire [7:0] _char_baseaddr_lut_T_7 = 3'h7 * 5'h10; // @[CharOutput.scala 110:60]
  wire [8:0] _char_baseaddr_lut_T_8 = 4'h8 * 5'h10; // @[CharOutput.scala 110:60]
  wire [8:0] _char_baseaddr_lut_T_9 = 4'h9 * 5'h10; // @[CharOutput.scala 110:60]
  wire [8:0] _char_baseaddr_lut_T_10 = 4'ha * 5'h10; // @[CharOutput.scala 110:60]
  wire [8:0] _char_baseaddr_lut_T_11 = 4'hb * 5'h10; // @[CharOutput.scala 110:60]
  wire [8:0] _char_baseaddr_lut_T_12 = 4'hc * 5'h10; // @[CharOutput.scala 110:60]
  wire [8:0] _char_baseaddr_lut_T_13 = 4'hd * 5'h10; // @[CharOutput.scala 110:60]
  wire [8:0] _char_baseaddr_lut_T_14 = 4'he * 5'h10; // @[CharOutput.scala 110:60]
  wire [8:0] _char_baseaddr_lut_T_15 = 4'hf * 5'h10; // @[CharOutput.scala 110:60]
  wire [9:0] _char_baseaddr_lut_T_16 = 5'h10 * 5'h10; // @[CharOutput.scala 110:60]
  wire [9:0] _char_baseaddr_lut_T_17 = 5'h11 * 5'h10; // @[CharOutput.scala 110:60]
  wire [9:0] _char_baseaddr_lut_T_18 = 5'h12 * 5'h10; // @[CharOutput.scala 110:60]
  wire [9:0] _char_baseaddr_lut_T_19 = 5'h13 * 5'h10; // @[CharOutput.scala 110:60]
  wire [9:0] _char_baseaddr_lut_T_20 = 5'h14 * 5'h10; // @[CharOutput.scala 110:60]
  wire [9:0] _char_baseaddr_lut_T_21 = 5'h15 * 5'h10; // @[CharOutput.scala 110:60]
  wire [9:0] _char_baseaddr_lut_T_22 = 5'h16 * 5'h10; // @[CharOutput.scala 110:60]
  wire [9:0] _char_baseaddr_lut_T_23 = 5'h17 * 5'h10; // @[CharOutput.scala 110:60]
  wire [9:0] _char_baseaddr_lut_T_24 = 5'h18 * 5'h10; // @[CharOutput.scala 110:60]
  wire [9:0] _char_baseaddr_lut_T_25 = 5'h19 * 5'h10; // @[CharOutput.scala 110:60]
  wire [9:0] _char_baseaddr_lut_T_26 = 5'h1a * 5'h10; // @[CharOutput.scala 110:60]
  wire [9:0] _char_baseaddr_lut_T_27 = 5'h1b * 5'h10; // @[CharOutput.scala 110:60]
  wire [9:0] _char_baseaddr_lut_T_28 = 5'h1c * 5'h10; // @[CharOutput.scala 110:60]
  wire [9:0] _char_baseaddr_lut_T_29 = 5'h1d * 5'h10; // @[CharOutput.scala 110:60]
  wire [9:0] _char_baseaddr_lut_T_30 = 5'h1e * 5'h10; // @[CharOutput.scala 110:60]
  wire [9:0] _char_baseaddr_lut_T_31 = 5'h1f * 5'h10; // @[CharOutput.scala 110:60]
  wire [10:0] _char_baseaddr_lut_T_32 = 6'h20 * 5'h10; // @[CharOutput.scala 110:60]
  wire [10:0] _char_baseaddr_lut_T_33 = 6'h21 * 5'h10; // @[CharOutput.scala 110:60]
  wire [10:0] _char_baseaddr_lut_T_34 = 6'h22 * 5'h10; // @[CharOutput.scala 110:60]
  wire [10:0] _char_baseaddr_lut_T_35 = 6'h23 * 5'h10; // @[CharOutput.scala 110:60]
  wire [10:0] _char_baseaddr_lut_T_36 = 6'h24 * 5'h10; // @[CharOutput.scala 110:60]
  wire [10:0] _char_baseaddr_lut_T_37 = 6'h25 * 5'h10; // @[CharOutput.scala 110:60]
  wire [10:0] _char_baseaddr_lut_T_38 = 6'h26 * 5'h10; // @[CharOutput.scala 110:60]
  wire [10:0] _char_baseaddr_lut_T_39 = 6'h27 * 5'h10; // @[CharOutput.scala 110:60]
  wire [10:0] _char_baseaddr_lut_T_40 = 6'h28 * 5'h10; // @[CharOutput.scala 110:60]
  wire [10:0] _char_baseaddr_lut_T_41 = 6'h29 * 5'h10; // @[CharOutput.scala 110:60]
  wire [10:0] _char_baseaddr_lut_T_42 = 6'h2a * 5'h10; // @[CharOutput.scala 110:60]
  wire [10:0] _char_baseaddr_lut_T_43 = 6'h2b * 5'h10; // @[CharOutput.scala 110:60]
  wire [10:0] _char_baseaddr_lut_T_44 = 6'h2c * 5'h10; // @[CharOutput.scala 110:60]
  wire [10:0] _char_baseaddr_lut_T_45 = 6'h2d * 5'h10; // @[CharOutput.scala 110:60]
  wire [10:0] _char_baseaddr_lut_T_46 = 6'h2e * 5'h10; // @[CharOutput.scala 110:60]
  wire [10:0] _char_baseaddr_lut_T_47 = 6'h2f * 5'h10; // @[CharOutput.scala 110:60]
  wire [10:0] _char_baseaddr_lut_T_48 = 6'h30 * 5'h10; // @[CharOutput.scala 110:60]
  wire [10:0] _char_baseaddr_lut_T_49 = 6'h31 * 5'h10; // @[CharOutput.scala 110:60]
  wire [10:0] _char_baseaddr_lut_T_50 = 6'h32 * 5'h10; // @[CharOutput.scala 110:60]
  wire [10:0] _char_baseaddr_lut_T_51 = 6'h33 * 5'h10; // @[CharOutput.scala 110:60]
  wire [10:0] _char_baseaddr_lut_T_52 = 6'h34 * 5'h10; // @[CharOutput.scala 110:60]
  wire [10:0] _char_baseaddr_lut_T_53 = 6'h35 * 5'h10; // @[CharOutput.scala 110:60]
  wire [10:0] _char_baseaddr_lut_T_54 = 6'h36 * 5'h10; // @[CharOutput.scala 110:60]
  wire [10:0] _char_baseaddr_lut_T_55 = 6'h37 * 5'h10; // @[CharOutput.scala 110:60]
  wire [10:0] _char_baseaddr_lut_T_56 = 6'h38 * 5'h10; // @[CharOutput.scala 110:60]
  wire [10:0] _char_baseaddr_lut_T_57 = 6'h39 * 5'h10; // @[CharOutput.scala 110:60]
  wire [10:0] _char_baseaddr_lut_T_58 = 6'h3a * 5'h10; // @[CharOutput.scala 110:60]
  wire [10:0] _char_baseaddr_lut_T_59 = 6'h3b * 5'h10; // @[CharOutput.scala 110:60]
  wire [10:0] _char_baseaddr_lut_T_60 = 6'h3c * 5'h10; // @[CharOutput.scala 110:60]
  wire [10:0] _char_baseaddr_lut_T_61 = 6'h3d * 5'h10; // @[CharOutput.scala 110:60]
  wire [10:0] _char_baseaddr_lut_T_62 = 6'h3e * 5'h10; // @[CharOutput.scala 110:60]
  wire [10:0] _char_baseaddr_lut_T_63 = 6'h3f * 5'h10; // @[CharOutput.scala 110:60]
  wire [11:0] _char_baseaddr_lut_T_64 = 7'h40 * 5'h10; // @[CharOutput.scala 110:60]
  wire [11:0] _char_baseaddr_lut_T_65 = 7'h41 * 5'h10; // @[CharOutput.scala 110:60]
  wire [11:0] _char_baseaddr_lut_T_66 = 7'h42 * 5'h10; // @[CharOutput.scala 110:60]
  wire [11:0] _char_baseaddr_lut_T_67 = 7'h43 * 5'h10; // @[CharOutput.scala 110:60]
  wire [11:0] _char_baseaddr_lut_T_68 = 7'h44 * 5'h10; // @[CharOutput.scala 110:60]
  wire [11:0] _char_baseaddr_lut_T_69 = 7'h45 * 5'h10; // @[CharOutput.scala 110:60]
  wire [11:0] _char_baseaddr_lut_T_70 = 7'h46 * 5'h10; // @[CharOutput.scala 110:60]
  wire [11:0] _char_baseaddr_lut_T_71 = 7'h47 * 5'h10; // @[CharOutput.scala 110:60]
  wire [11:0] _char_baseaddr_lut_T_72 = 7'h48 * 5'h10; // @[CharOutput.scala 110:60]
  wire [11:0] _char_baseaddr_lut_T_73 = 7'h49 * 5'h10; // @[CharOutput.scala 110:60]
  wire [11:0] _char_baseaddr_lut_T_74 = 7'h4a * 5'h10; // @[CharOutput.scala 110:60]
  wire [11:0] _char_baseaddr_lut_T_75 = 7'h4b * 5'h10; // @[CharOutput.scala 110:60]
  wire [11:0] _char_baseaddr_lut_T_76 = 7'h4c * 5'h10; // @[CharOutput.scala 110:60]
  wire [11:0] _char_baseaddr_lut_T_77 = 7'h4d * 5'h10; // @[CharOutput.scala 110:60]
  wire [11:0] _char_baseaddr_lut_T_78 = 7'h4e * 5'h10; // @[CharOutput.scala 110:60]
  wire [11:0] _char_baseaddr_lut_T_79 = 7'h4f * 5'h10; // @[CharOutput.scala 110:60]
  wire [11:0] _char_baseaddr_lut_T_80 = 7'h50 * 5'h10; // @[CharOutput.scala 110:60]
  wire [11:0] _char_baseaddr_lut_T_81 = 7'h51 * 5'h10; // @[CharOutput.scala 110:60]
  wire [11:0] _char_baseaddr_lut_T_82 = 7'h52 * 5'h10; // @[CharOutput.scala 110:60]
  wire [11:0] _char_baseaddr_lut_T_83 = 7'h53 * 5'h10; // @[CharOutput.scala 110:60]
  wire [11:0] _char_baseaddr_lut_T_84 = 7'h54 * 5'h10; // @[CharOutput.scala 110:60]
  wire [11:0] _char_baseaddr_lut_T_85 = 7'h55 * 5'h10; // @[CharOutput.scala 110:60]
  wire [11:0] _char_baseaddr_lut_T_86 = 7'h56 * 5'h10; // @[CharOutput.scala 110:60]
  wire [11:0] _char_baseaddr_lut_T_87 = 7'h57 * 5'h10; // @[CharOutput.scala 110:60]
  wire [11:0] _char_baseaddr_lut_T_88 = 7'h58 * 5'h10; // @[CharOutput.scala 110:60]
  wire [11:0] _char_baseaddr_lut_T_89 = 7'h59 * 5'h10; // @[CharOutput.scala 110:60]
  wire [11:0] _char_baseaddr_lut_T_90 = 7'h5a * 5'h10; // @[CharOutput.scala 110:60]
  wire [11:0] _char_baseaddr_lut_T_91 = 7'h5b * 5'h10; // @[CharOutput.scala 110:60]
  wire [11:0] _char_baseaddr_lut_T_92 = 7'h5c * 5'h10; // @[CharOutput.scala 110:60]
  wire [11:0] _char_baseaddr_lut_T_93 = 7'h5d * 5'h10; // @[CharOutput.scala 110:60]
  wire [11:0] _char_baseaddr_lut_T_94 = 7'h5e * 5'h10; // @[CharOutput.scala 110:60]
  wire [11:0] _char_baseaddr_lut_T_95 = 7'h5f * 5'h10; // @[CharOutput.scala 110:60]
  wire [11:0] _char_baseaddr_lut_T_96 = 7'h60 * 5'h10; // @[CharOutput.scala 110:60]
  wire [11:0] _char_baseaddr_lut_T_97 = 7'h61 * 5'h10; // @[CharOutput.scala 110:60]
  wire [11:0] _char_baseaddr_lut_T_98 = 7'h62 * 5'h10; // @[CharOutput.scala 110:60]
  wire [11:0] _char_baseaddr_lut_T_99 = 7'h63 * 5'h10; // @[CharOutput.scala 110:60]
  wire [11:0] _char_baseaddr_lut_T_100 = 7'h64 * 5'h10; // @[CharOutput.scala 110:60]
  wire [11:0] _char_baseaddr_lut_T_101 = 7'h65 * 5'h10; // @[CharOutput.scala 110:60]
  wire [11:0] _char_baseaddr_lut_T_102 = 7'h66 * 5'h10; // @[CharOutput.scala 110:60]
  wire [11:0] _char_baseaddr_lut_T_103 = 7'h67 * 5'h10; // @[CharOutput.scala 110:60]
  wire [11:0] _char_baseaddr_lut_T_104 = 7'h68 * 5'h10; // @[CharOutput.scala 110:60]
  wire [11:0] _char_baseaddr_lut_T_105 = 7'h69 * 5'h10; // @[CharOutput.scala 110:60]
  wire [11:0] _char_baseaddr_lut_T_106 = 7'h6a * 5'h10; // @[CharOutput.scala 110:60]
  wire [11:0] _char_baseaddr_lut_T_107 = 7'h6b * 5'h10; // @[CharOutput.scala 110:60]
  wire [11:0] _char_baseaddr_lut_T_108 = 7'h6c * 5'h10; // @[CharOutput.scala 110:60]
  wire [11:0] _char_baseaddr_lut_T_109 = 7'h6d * 5'h10; // @[CharOutput.scala 110:60]
  wire [11:0] _char_baseaddr_lut_T_110 = 7'h6e * 5'h10; // @[CharOutput.scala 110:60]
  wire [11:0] _char_baseaddr_lut_T_111 = 7'h6f * 5'h10; // @[CharOutput.scala 110:60]
  wire [11:0] _char_baseaddr_lut_T_112 = 7'h70 * 5'h10; // @[CharOutput.scala 110:60]
  wire [11:0] _char_baseaddr_lut_T_113 = 7'h71 * 5'h10; // @[CharOutput.scala 110:60]
  wire [11:0] _char_baseaddr_lut_T_114 = 7'h72 * 5'h10; // @[CharOutput.scala 110:60]
  wire [11:0] _char_baseaddr_lut_T_115 = 7'h73 * 5'h10; // @[CharOutput.scala 110:60]
  wire [11:0] _char_baseaddr_lut_T_116 = 7'h74 * 5'h10; // @[CharOutput.scala 110:60]
  wire [11:0] _char_baseaddr_lut_T_117 = 7'h75 * 5'h10; // @[CharOutput.scala 110:60]
  wire [11:0] _char_baseaddr_lut_T_118 = 7'h76 * 5'h10; // @[CharOutput.scala 110:60]
  wire [11:0] _char_baseaddr_lut_T_119 = 7'h77 * 5'h10; // @[CharOutput.scala 110:60]
  wire [11:0] _char_baseaddr_lut_T_120 = 7'h78 * 5'h10; // @[CharOutput.scala 110:60]
  wire [11:0] _char_baseaddr_lut_T_121 = 7'h79 * 5'h10; // @[CharOutput.scala 110:60]
  wire [11:0] _char_baseaddr_lut_T_122 = 7'h7a * 5'h10; // @[CharOutput.scala 110:60]
  wire [11:0] _char_baseaddr_lut_T_123 = 7'h7b * 5'h10; // @[CharOutput.scala 110:60]
  wire [11:0] _char_baseaddr_lut_T_124 = 7'h7c * 5'h10; // @[CharOutput.scala 110:60]
  wire [11:0] _char_baseaddr_lut_T_125 = 7'h7d * 5'h10; // @[CharOutput.scala 110:60]
  wire [11:0] _char_baseaddr_lut_T_126 = 7'h7e * 5'h10; // @[CharOutput.scala 110:60]
  wire [11:0] _char_baseaddr_lut_T_127 = 7'h7f * 5'h10; // @[CharOutput.scala 110:60]
  wire [12:0] char_baseaddr_lut_128 = 8'h80 * 5'h10; // @[CharOutput.scala 110:60]
  wire [12:0] char_baseaddr_lut_129 = 8'h81 * 5'h10; // @[CharOutput.scala 110:60]
  wire [12:0] char_baseaddr_lut_130 = 8'h82 * 5'h10; // @[CharOutput.scala 110:60]
  wire [12:0] char_baseaddr_lut_131 = 8'h83 * 5'h10; // @[CharOutput.scala 110:60]
  wire [12:0] char_baseaddr_lut_132 = 8'h84 * 5'h10; // @[CharOutput.scala 110:60]
  wire [12:0] char_baseaddr_lut_133 = 8'h85 * 5'h10; // @[CharOutput.scala 110:60]
  wire [12:0] char_baseaddr_lut_134 = 8'h86 * 5'h10; // @[CharOutput.scala 110:60]
  wire [12:0] char_baseaddr_lut_135 = 8'h87 * 5'h10; // @[CharOutput.scala 110:60]
  wire [12:0] char_baseaddr_lut_136 = 8'h88 * 5'h10; // @[CharOutput.scala 110:60]
  wire [12:0] char_baseaddr_lut_137 = 8'h89 * 5'h10; // @[CharOutput.scala 110:60]
  wire [12:0] char_baseaddr_lut_138 = 8'h8a * 5'h10; // @[CharOutput.scala 110:60]
  wire [12:0] char_baseaddr_lut_139 = 8'h8b * 5'h10; // @[CharOutput.scala 110:60]
  wire [12:0] char_baseaddr_lut_140 = 8'h8c * 5'h10; // @[CharOutput.scala 110:60]
  wire [12:0] char_baseaddr_lut_141 = 8'h8d * 5'h10; // @[CharOutput.scala 110:60]
  wire [12:0] char_baseaddr_lut_142 = 8'h8e * 5'h10; // @[CharOutput.scala 110:60]
  wire [12:0] char_baseaddr_lut_143 = 8'h8f * 5'h10; // @[CharOutput.scala 110:60]
  wire [12:0] char_baseaddr_lut_144 = 8'h90 * 5'h10; // @[CharOutput.scala 110:60]
  wire [12:0] char_baseaddr_lut_145 = 8'h91 * 5'h10; // @[CharOutput.scala 110:60]
  wire [12:0] char_baseaddr_lut_146 = 8'h92 * 5'h10; // @[CharOutput.scala 110:60]
  wire [12:0] char_baseaddr_lut_147 = 8'h93 * 5'h10; // @[CharOutput.scala 110:60]
  wire [12:0] char_baseaddr_lut_148 = 8'h94 * 5'h10; // @[CharOutput.scala 110:60]
  wire [12:0] char_baseaddr_lut_149 = 8'h95 * 5'h10; // @[CharOutput.scala 110:60]
  wire [12:0] char_baseaddr_lut_150 = 8'h96 * 5'h10; // @[CharOutput.scala 110:60]
  wire [12:0] char_baseaddr_lut_151 = 8'h97 * 5'h10; // @[CharOutput.scala 110:60]
  wire [12:0] char_baseaddr_lut_152 = 8'h98 * 5'h10; // @[CharOutput.scala 110:60]
  wire [12:0] char_baseaddr_lut_153 = 8'h99 * 5'h10; // @[CharOutput.scala 110:60]
  wire [12:0] char_baseaddr_lut_154 = 8'h9a * 5'h10; // @[CharOutput.scala 110:60]
  wire [12:0] char_baseaddr_lut_155 = 8'h9b * 5'h10; // @[CharOutput.scala 110:60]
  wire [12:0] char_baseaddr_lut_156 = 8'h9c * 5'h10; // @[CharOutput.scala 110:60]
  wire [12:0] char_baseaddr_lut_157 = 8'h9d * 5'h10; // @[CharOutput.scala 110:60]
  wire [12:0] char_baseaddr_lut_158 = 8'h9e * 5'h10; // @[CharOutput.scala 110:60]
  wire [12:0] char_baseaddr_lut_159 = 8'h9f * 5'h10; // @[CharOutput.scala 110:60]
  wire [12:0] char_baseaddr_lut_160 = 8'ha0 * 5'h10; // @[CharOutput.scala 110:60]
  wire [12:0] char_baseaddr_lut_161 = 8'ha1 * 5'h10; // @[CharOutput.scala 110:60]
  wire [12:0] char_baseaddr_lut_162 = 8'ha2 * 5'h10; // @[CharOutput.scala 110:60]
  wire [12:0] char_baseaddr_lut_163 = 8'ha3 * 5'h10; // @[CharOutput.scala 110:60]
  wire [12:0] char_baseaddr_lut_164 = 8'ha4 * 5'h10; // @[CharOutput.scala 110:60]
  wire [12:0] char_baseaddr_lut_165 = 8'ha5 * 5'h10; // @[CharOutput.scala 110:60]
  wire [12:0] char_baseaddr_lut_166 = 8'ha6 * 5'h10; // @[CharOutput.scala 110:60]
  wire [12:0] char_baseaddr_lut_167 = 8'ha7 * 5'h10; // @[CharOutput.scala 110:60]
  wire [12:0] char_baseaddr_lut_168 = 8'ha8 * 5'h10; // @[CharOutput.scala 110:60]
  wire [12:0] char_baseaddr_lut_169 = 8'ha9 * 5'h10; // @[CharOutput.scala 110:60]
  wire [12:0] char_baseaddr_lut_170 = 8'haa * 5'h10; // @[CharOutput.scala 110:60]
  wire [12:0] char_baseaddr_lut_171 = 8'hab * 5'h10; // @[CharOutput.scala 110:60]
  wire [12:0] char_baseaddr_lut_172 = 8'hac * 5'h10; // @[CharOutput.scala 110:60]
  wire [12:0] char_baseaddr_lut_173 = 8'had * 5'h10; // @[CharOutput.scala 110:60]
  wire [12:0] char_baseaddr_lut_174 = 8'hae * 5'h10; // @[CharOutput.scala 110:60]
  wire [12:0] char_baseaddr_lut_175 = 8'haf * 5'h10; // @[CharOutput.scala 110:60]
  wire [12:0] char_baseaddr_lut_176 = 8'hb0 * 5'h10; // @[CharOutput.scala 110:60]
  wire [12:0] char_baseaddr_lut_177 = 8'hb1 * 5'h10; // @[CharOutput.scala 110:60]
  wire [12:0] char_baseaddr_lut_178 = 8'hb2 * 5'h10; // @[CharOutput.scala 110:60]
  wire [12:0] char_baseaddr_lut_179 = 8'hb3 * 5'h10; // @[CharOutput.scala 110:60]
  wire [12:0] char_baseaddr_lut_180 = 8'hb4 * 5'h10; // @[CharOutput.scala 110:60]
  wire [12:0] char_baseaddr_lut_181 = 8'hb5 * 5'h10; // @[CharOutput.scala 110:60]
  wire [12:0] char_baseaddr_lut_182 = 8'hb6 * 5'h10; // @[CharOutput.scala 110:60]
  wire [12:0] char_baseaddr_lut_183 = 8'hb7 * 5'h10; // @[CharOutput.scala 110:60]
  wire [12:0] char_baseaddr_lut_184 = 8'hb8 * 5'h10; // @[CharOutput.scala 110:60]
  wire [12:0] char_baseaddr_lut_185 = 8'hb9 * 5'h10; // @[CharOutput.scala 110:60]
  wire [12:0] char_baseaddr_lut_186 = 8'hba * 5'h10; // @[CharOutput.scala 110:60]
  wire [12:0] char_baseaddr_lut_187 = 8'hbb * 5'h10; // @[CharOutput.scala 110:60]
  wire [12:0] char_baseaddr_lut_188 = 8'hbc * 5'h10; // @[CharOutput.scala 110:60]
  wire [12:0] char_baseaddr_lut_189 = 8'hbd * 5'h10; // @[CharOutput.scala 110:60]
  wire [12:0] char_baseaddr_lut_190 = 8'hbe * 5'h10; // @[CharOutput.scala 110:60]
  wire [12:0] char_baseaddr_lut_191 = 8'hbf * 5'h10; // @[CharOutput.scala 110:60]
  wire [12:0] char_baseaddr_lut_192 = 8'hc0 * 5'h10; // @[CharOutput.scala 110:60]
  wire [12:0] char_baseaddr_lut_193 = 8'hc1 * 5'h10; // @[CharOutput.scala 110:60]
  wire [12:0] char_baseaddr_lut_194 = 8'hc2 * 5'h10; // @[CharOutput.scala 110:60]
  wire [12:0] char_baseaddr_lut_195 = 8'hc3 * 5'h10; // @[CharOutput.scala 110:60]
  wire [12:0] char_baseaddr_lut_196 = 8'hc4 * 5'h10; // @[CharOutput.scala 110:60]
  wire [12:0] char_baseaddr_lut_197 = 8'hc5 * 5'h10; // @[CharOutput.scala 110:60]
  wire [12:0] char_baseaddr_lut_198 = 8'hc6 * 5'h10; // @[CharOutput.scala 110:60]
  wire [12:0] char_baseaddr_lut_199 = 8'hc7 * 5'h10; // @[CharOutput.scala 110:60]
  wire [12:0] char_baseaddr_lut_200 = 8'hc8 * 5'h10; // @[CharOutput.scala 110:60]
  wire [12:0] char_baseaddr_lut_201 = 8'hc9 * 5'h10; // @[CharOutput.scala 110:60]
  wire [12:0] char_baseaddr_lut_202 = 8'hca * 5'h10; // @[CharOutput.scala 110:60]
  wire [12:0] char_baseaddr_lut_203 = 8'hcb * 5'h10; // @[CharOutput.scala 110:60]
  wire [12:0] char_baseaddr_lut_204 = 8'hcc * 5'h10; // @[CharOutput.scala 110:60]
  wire [12:0] char_baseaddr_lut_205 = 8'hcd * 5'h10; // @[CharOutput.scala 110:60]
  wire [12:0] char_baseaddr_lut_206 = 8'hce * 5'h10; // @[CharOutput.scala 110:60]
  wire [12:0] char_baseaddr_lut_207 = 8'hcf * 5'h10; // @[CharOutput.scala 110:60]
  wire [12:0] char_baseaddr_lut_208 = 8'hd0 * 5'h10; // @[CharOutput.scala 110:60]
  wire [12:0] char_baseaddr_lut_209 = 8'hd1 * 5'h10; // @[CharOutput.scala 110:60]
  wire [12:0] char_baseaddr_lut_210 = 8'hd2 * 5'h10; // @[CharOutput.scala 110:60]
  wire [12:0] char_baseaddr_lut_211 = 8'hd3 * 5'h10; // @[CharOutput.scala 110:60]
  wire [12:0] char_baseaddr_lut_212 = 8'hd4 * 5'h10; // @[CharOutput.scala 110:60]
  wire [12:0] char_baseaddr_lut_213 = 8'hd5 * 5'h10; // @[CharOutput.scala 110:60]
  wire [12:0] char_baseaddr_lut_214 = 8'hd6 * 5'h10; // @[CharOutput.scala 110:60]
  wire [12:0] char_baseaddr_lut_215 = 8'hd7 * 5'h10; // @[CharOutput.scala 110:60]
  wire [12:0] char_baseaddr_lut_216 = 8'hd8 * 5'h10; // @[CharOutput.scala 110:60]
  wire [12:0] char_baseaddr_lut_217 = 8'hd9 * 5'h10; // @[CharOutput.scala 110:60]
  wire [12:0] char_baseaddr_lut_218 = 8'hda * 5'h10; // @[CharOutput.scala 110:60]
  wire [12:0] char_baseaddr_lut_219 = 8'hdb * 5'h10; // @[CharOutput.scala 110:60]
  wire [12:0] char_baseaddr_lut_220 = 8'hdc * 5'h10; // @[CharOutput.scala 110:60]
  wire [12:0] char_baseaddr_lut_221 = 8'hdd * 5'h10; // @[CharOutput.scala 110:60]
  wire [12:0] char_baseaddr_lut_222 = 8'hde * 5'h10; // @[CharOutput.scala 110:60]
  wire [12:0] char_baseaddr_lut_223 = 8'hdf * 5'h10; // @[CharOutput.scala 110:60]
  wire [12:0] char_baseaddr_lut_224 = 8'he0 * 5'h10; // @[CharOutput.scala 110:60]
  wire [12:0] char_baseaddr_lut_225 = 8'he1 * 5'h10; // @[CharOutput.scala 110:60]
  wire [12:0] char_baseaddr_lut_226 = 8'he2 * 5'h10; // @[CharOutput.scala 110:60]
  wire [12:0] char_baseaddr_lut_227 = 8'he3 * 5'h10; // @[CharOutput.scala 110:60]
  wire [12:0] char_baseaddr_lut_228 = 8'he4 * 5'h10; // @[CharOutput.scala 110:60]
  wire [12:0] char_baseaddr_lut_229 = 8'he5 * 5'h10; // @[CharOutput.scala 110:60]
  wire [12:0] char_baseaddr_lut_230 = 8'he6 * 5'h10; // @[CharOutput.scala 110:60]
  wire [12:0] char_baseaddr_lut_231 = 8'he7 * 5'h10; // @[CharOutput.scala 110:60]
  wire [12:0] char_baseaddr_lut_232 = 8'he8 * 5'h10; // @[CharOutput.scala 110:60]
  wire [12:0] char_baseaddr_lut_233 = 8'he9 * 5'h10; // @[CharOutput.scala 110:60]
  wire [12:0] char_baseaddr_lut_234 = 8'hea * 5'h10; // @[CharOutput.scala 110:60]
  wire [12:0] char_baseaddr_lut_235 = 8'heb * 5'h10; // @[CharOutput.scala 110:60]
  wire [12:0] char_baseaddr_lut_236 = 8'hec * 5'h10; // @[CharOutput.scala 110:60]
  wire [12:0] char_baseaddr_lut_237 = 8'hed * 5'h10; // @[CharOutput.scala 110:60]
  wire [12:0] char_baseaddr_lut_238 = 8'hee * 5'h10; // @[CharOutput.scala 110:60]
  wire [12:0] char_baseaddr_lut_239 = 8'hef * 5'h10; // @[CharOutput.scala 110:60]
  wire [12:0] char_baseaddr_lut_240 = 8'hf0 * 5'h10; // @[CharOutput.scala 110:60]
  wire [12:0] char_baseaddr_lut_241 = 8'hf1 * 5'h10; // @[CharOutput.scala 110:60]
  wire [12:0] char_baseaddr_lut_242 = 8'hf2 * 5'h10; // @[CharOutput.scala 110:60]
  wire [12:0] char_baseaddr_lut_243 = 8'hf3 * 5'h10; // @[CharOutput.scala 110:60]
  wire [12:0] char_baseaddr_lut_244 = 8'hf4 * 5'h10; // @[CharOutput.scala 110:60]
  wire [12:0] char_baseaddr_lut_245 = 8'hf5 * 5'h10; // @[CharOutput.scala 110:60]
  wire [12:0] char_baseaddr_lut_246 = 8'hf6 * 5'h10; // @[CharOutput.scala 110:60]
  wire [12:0] char_baseaddr_lut_247 = 8'hf7 * 5'h10; // @[CharOutput.scala 110:60]
  wire [12:0] char_baseaddr_lut_248 = 8'hf8 * 5'h10; // @[CharOutput.scala 110:60]
  wire [12:0] char_baseaddr_lut_249 = 8'hf9 * 5'h10; // @[CharOutput.scala 110:60]
  wire [12:0] char_baseaddr_lut_250 = 8'hfa * 5'h10; // @[CharOutput.scala 110:60]
  wire [12:0] char_baseaddr_lut_251 = 8'hfb * 5'h10; // @[CharOutput.scala 110:60]
  wire [12:0] char_baseaddr_lut_252 = 8'hfc * 5'h10; // @[CharOutput.scala 110:60]
  wire [12:0] char_baseaddr_lut_253 = 8'hfd * 5'h10; // @[CharOutput.scala 110:60]
  wire [12:0] char_baseaddr_lut_254 = 8'hfe * 5'h10; // @[CharOutput.scala 110:60]
  wire [12:0] char_baseaddr_lut_255 = 8'hff * 5'h10; // @[CharOutput.scala 110:60]
  wire [4:0] _GEN_1112 = 3'h1 == obj_choose ? io_class_voc_1 : io_class_voc_0; // @[CharOutput.scala 115:{23,23}]
  wire [4:0] _GEN_1113 = 3'h2 == obj_choose ? io_class_voc_2 : _GEN_1112; // @[CharOutput.scala 115:{23,23}]
  wire [4:0] _GEN_1114 = 3'h3 == obj_choose ? io_class_voc_3 : _GEN_1113; // @[CharOutput.scala 115:{23,23}]
  wire [4:0] _GEN_1115 = 3'h4 == obj_choose ? io_class_voc_4 : _GEN_1114; // @[CharOutput.scala 115:{23,23}]
  wire [7:0] _GEN_1117 = 5'h1 == _GEN_1115 ? 8'h62 : 8'h41; // @[CharOutput.scala 115:{23,23}]
  wire [7:0] _GEN_1118 = 5'h2 == _GEN_1115 ? 8'h62 : _GEN_1117; // @[CharOutput.scala 115:{23,23}]
  wire [7:0] _GEN_1119 = 5'h3 == _GEN_1115 ? 8'h62 : _GEN_1118; // @[CharOutput.scala 115:{23,23}]
  wire [7:0] _GEN_1120 = 5'h4 == _GEN_1115 ? 8'h62 : _GEN_1119; // @[CharOutput.scala 115:{23,23}]
  wire [7:0] _GEN_1121 = 5'h5 == _GEN_1115 ? 8'h62 : _GEN_1120; // @[CharOutput.scala 115:{23,23}]
  wire [7:0] _GEN_1122 = 5'h6 == _GEN_1115 ? 8'h63 : _GEN_1121; // @[CharOutput.scala 115:{23,23}]
  wire [7:0] _GEN_1123 = 5'h7 == _GEN_1115 ? 8'h63 : _GEN_1122; // @[CharOutput.scala 115:{23,23}]
  wire [7:0] _GEN_1124 = 5'h8 == _GEN_1115 ? 8'h63 : _GEN_1123; // @[CharOutput.scala 115:{23,23}]
  wire [7:0] _GEN_1125 = 5'h9 == _GEN_1115 ? 8'h63 : _GEN_1124; // @[CharOutput.scala 115:{23,23}]
  wire [7:0] _GEN_1126 = 5'ha == _GEN_1115 ? 8'h64 : _GEN_1125; // @[CharOutput.scala 115:{23,23}]
  wire [7:0] _GEN_1127 = 5'hb == _GEN_1115 ? 8'h64 : _GEN_1126; // @[CharOutput.scala 115:{23,23}]
  wire [7:0] _GEN_1128 = 5'hc == _GEN_1115 ? 8'h68 : _GEN_1127; // @[CharOutput.scala 115:{23,23}]
  wire [7:0] _GEN_1129 = 5'hd == _GEN_1115 ? 8'h6d : _GEN_1128; // @[CharOutput.scala 115:{23,23}]
  wire [7:0] _GEN_1130 = 5'he == _GEN_1115 ? 8'h70 : _GEN_1129; // @[CharOutput.scala 115:{23,23}]
  wire [7:0] _GEN_1131 = 5'hf == _GEN_1115 ? 8'h70 : _GEN_1130; // @[CharOutput.scala 115:{23,23}]
  wire [7:0] _GEN_1132 = 5'h10 == _GEN_1115 ? 8'h73 : _GEN_1131; // @[CharOutput.scala 115:{23,23}]
  wire [7:0] _GEN_1133 = 5'h11 == _GEN_1115 ? 8'h73 : _GEN_1132; // @[CharOutput.scala 115:{23,23}]
  wire [7:0] _GEN_1134 = 5'h12 == _GEN_1115 ? 8'h74 : _GEN_1133; // @[CharOutput.scala 115:{23,23}]
  wire [7:0] current_ascii_array_0 = 5'h13 == _GEN_1115 ? 8'h74 : _GEN_1134; // @[CharOutput.scala 115:{23,23}]
  wire [7:0] _GEN_1137 = 5'h1 == _GEN_1115 ? 8'h69 : 8'h65; // @[CharOutput.scala 115:{23,23}]
  wire [7:0] _GEN_1138 = 5'h2 == _GEN_1115 ? 8'h69 : _GEN_1137; // @[CharOutput.scala 115:{23,23}]
  wire [7:0] _GEN_1139 = 5'h3 == _GEN_1115 ? 8'h6f : _GEN_1138; // @[CharOutput.scala 115:{23,23}]
  wire [7:0] _GEN_1140 = 5'h4 == _GEN_1115 ? 8'h6f : _GEN_1139; // @[CharOutput.scala 115:{23,23}]
  wire [7:0] _GEN_1141 = 5'h5 == _GEN_1115 ? 8'h75 : _GEN_1140; // @[CharOutput.scala 115:{23,23}]
  wire [7:0] _GEN_1142 = 5'h6 == _GEN_1115 ? 8'h61 : _GEN_1141; // @[CharOutput.scala 115:{23,23}]
  wire [7:0] _GEN_1143 = 5'h7 == _GEN_1115 ? 8'h61 : _GEN_1142; // @[CharOutput.scala 115:{23,23}]
  wire [7:0] _GEN_1144 = 5'h8 == _GEN_1115 ? 8'h68 : _GEN_1143; // @[CharOutput.scala 115:{23,23}]
  wire [7:0] _GEN_1145 = 5'h9 == _GEN_1115 ? 8'h6f : _GEN_1144; // @[CharOutput.scala 115:{23,23}]
  wire [7:0] _GEN_1146 = 5'ha == _GEN_1115 ? 8'h69 : _GEN_1145; // @[CharOutput.scala 115:{23,23}]
  wire [7:0] _GEN_1147 = 5'hb == _GEN_1115 ? 8'h6f : _GEN_1146; // @[CharOutput.scala 115:{23,23}]
  wire [7:0] _GEN_1148 = 5'hc == _GEN_1115 ? 8'h6f : _GEN_1147; // @[CharOutput.scala 115:{23,23}]
  wire [7:0] _GEN_1149 = 5'hd == _GEN_1115 ? 8'h6f : _GEN_1148; // @[CharOutput.scala 115:{23,23}]
  wire [7:0] _GEN_1150 = 5'he == _GEN_1115 ? 8'h65 : _GEN_1149; // @[CharOutput.scala 115:{23,23}]
  wire [7:0] _GEN_1151 = 5'hf == _GEN_1115 ? 8'h6f : _GEN_1150; // @[CharOutput.scala 115:{23,23}]
  wire [7:0] _GEN_1152 = 5'h10 == _GEN_1115 ? 8'h68 : _GEN_1151; // @[CharOutput.scala 115:{23,23}]
  wire [7:0] _GEN_1153 = 5'h11 == _GEN_1115 ? 8'h6f : _GEN_1152; // @[CharOutput.scala 115:{23,23}]
  wire [7:0] _GEN_1154 = 5'h12 == _GEN_1115 ? 8'h72 : _GEN_1153; // @[CharOutput.scala 115:{23,23}]
  wire [7:0] current_ascii_array_1 = 5'h13 == _GEN_1115 ? 8'h76 : _GEN_1154; // @[CharOutput.scala 115:{23,23}]
  wire [7:0] _GEN_1157 = 5'h1 == _GEN_1115 ? 8'h63 : 8'h72; // @[CharOutput.scala 115:{23,23}]
  wire [7:0] _GEN_1158 = 5'h2 == _GEN_1115 ? 8'h72 : _GEN_1157; // @[CharOutput.scala 115:{23,23}]
  wire [7:0] _GEN_1159 = 5'h3 == _GEN_1115 ? 8'h61 : _GEN_1158; // @[CharOutput.scala 115:{23,23}]
  wire [7:0] _GEN_1160 = 5'h4 == _GEN_1115 ? 8'h74 : _GEN_1159; // @[CharOutput.scala 115:{23,23}]
  wire [7:0] _GEN_1161 = 5'h5 == _GEN_1115 ? 8'h73 : _GEN_1160; // @[CharOutput.scala 115:{23,23}]
  wire [7:0] _GEN_1162 = 5'h6 == _GEN_1115 ? 8'h72 : _GEN_1161; // @[CharOutput.scala 115:{23,23}]
  wire [7:0] _GEN_1163 = 5'h7 == _GEN_1115 ? 8'h74 : _GEN_1162; // @[CharOutput.scala 115:{23,23}]
  wire [7:0] _GEN_1164 = 5'h8 == _GEN_1115 ? 8'h61 : _GEN_1163; // @[CharOutput.scala 115:{23,23}]
  wire [7:0] _GEN_1165 = 5'h9 == _GEN_1115 ? 8'h77 : _GEN_1164; // @[CharOutput.scala 115:{23,23}]
  wire [7:0] _GEN_1166 = 5'ha == _GEN_1115 ? 8'h6e : _GEN_1165; // @[CharOutput.scala 115:{23,23}]
  wire [7:0] _GEN_1167 = 5'hb == _GEN_1115 ? 8'h67 : _GEN_1166; // @[CharOutput.scala 115:{23,23}]
  wire [7:0] _GEN_1168 = 5'hc == _GEN_1115 ? 8'h72 : _GEN_1167; // @[CharOutput.scala 115:{23,23}]
  wire [7:0] _GEN_1169 = 5'hd == _GEN_1115 ? 8'h74 : _GEN_1168; // @[CharOutput.scala 115:{23,23}]
  wire [7:0] _GEN_1170 = 5'he == _GEN_1115 ? 8'h72 : _GEN_1169; // @[CharOutput.scala 115:{23,23}]
  wire [7:0] _GEN_1171 = 5'hf == _GEN_1115 ? 8'h74 : _GEN_1170; // @[CharOutput.scala 115:{23,23}]
  wire [7:0] _GEN_1172 = 5'h10 == _GEN_1115 ? 8'h65 : _GEN_1171; // @[CharOutput.scala 115:{23,23}]
  wire [7:0] _GEN_1173 = 5'h11 == _GEN_1115 ? 8'h66 : _GEN_1172; // @[CharOutput.scala 115:{23,23}]
  wire [7:0] _GEN_1174 = 5'h12 == _GEN_1115 ? 8'h61 : _GEN_1173; // @[CharOutput.scala 115:{23,23}]
  wire [7:0] current_ascii_array_2 = 5'h13 == _GEN_1115 ? 8'h6d : _GEN_1174; // @[CharOutput.scala 115:{23,23}]
  wire [7:0] _GEN_1177 = 5'h1 == _GEN_1115 ? 8'h79 : 8'h6f; // @[CharOutput.scala 115:{23,23}]
  wire [7:0] _GEN_1178 = 5'h2 == _GEN_1115 ? 8'h64 : _GEN_1177; // @[CharOutput.scala 115:{23,23}]
  wire [7:0] _GEN_1179 = 5'h3 == _GEN_1115 ? 8'h74 : _GEN_1178; // @[CharOutput.scala 115:{23,23}]
  wire [7:0] _GEN_1180 = 5'h4 == _GEN_1115 ? 8'h74 : _GEN_1179; // @[CharOutput.scala 115:{23,23}]
  wire [7:0] _GEN_1181 = 5'h5 == _GEN_1115 ? 8'h0 : _GEN_1180; // @[CharOutput.scala 115:{23,23}]
  wire [7:0] _GEN_1182 = 5'h6 == _GEN_1115 ? 8'h0 : _GEN_1181; // @[CharOutput.scala 115:{23,23}]
  wire [7:0] _GEN_1183 = 5'h7 == _GEN_1115 ? 8'h0 : _GEN_1182; // @[CharOutput.scala 115:{23,23}]
  wire [7:0] _GEN_1184 = 5'h8 == _GEN_1115 ? 8'h69 : _GEN_1183; // @[CharOutput.scala 115:{23,23}]
  wire [7:0] _GEN_1185 = 5'h9 == _GEN_1115 ? 8'h0 : _GEN_1184; // @[CharOutput.scala 115:{23,23}]
  wire [7:0] _GEN_1186 = 5'ha == _GEN_1115 ? 8'h69 : _GEN_1185; // @[CharOutput.scala 115:{23,23}]
  wire [7:0] _GEN_1187 = 5'hb == _GEN_1115 ? 8'h0 : _GEN_1186; // @[CharOutput.scala 115:{23,23}]
  wire [7:0] _GEN_1188 = 5'hc == _GEN_1115 ? 8'h73 : _GEN_1187; // @[CharOutput.scala 115:{23,23}]
  wire [7:0] _GEN_1189 = 5'hd == _GEN_1115 ? 8'h6f : _GEN_1188; // @[CharOutput.scala 115:{23,23}]
  wire [7:0] _GEN_1190 = 5'he == _GEN_1115 ? 8'h73 : _GEN_1189; // @[CharOutput.scala 115:{23,23}]
  wire [7:0] _GEN_1191 = 5'hf == _GEN_1115 ? 8'h74 : _GEN_1190; // @[CharOutput.scala 115:{23,23}]
  wire [7:0] _GEN_1192 = 5'h10 == _GEN_1115 ? 8'h65 : _GEN_1191; // @[CharOutput.scala 115:{23,23}]
  wire [7:0] _GEN_1193 = 5'h11 == _GEN_1115 ? 8'h61 : _GEN_1192; // @[CharOutput.scala 115:{23,23}]
  wire [7:0] _GEN_1194 = 5'h12 == _GEN_1115 ? 8'h69 : _GEN_1193; // @[CharOutput.scala 115:{23,23}]
  wire [7:0] current_ascii_array_3 = 5'h13 == _GEN_1115 ? 8'h6f : _GEN_1194; // @[CharOutput.scala 115:{23,23}]
  wire [7:0] _GEN_1197 = 5'h1 == _GEN_1115 ? 8'h63 : 8'h70; // @[CharOutput.scala 115:{23,23}]
  wire [7:0] _GEN_1198 = 5'h2 == _GEN_1115 ? 8'h0 : _GEN_1197; // @[CharOutput.scala 115:{23,23}]
  wire [7:0] _GEN_1199 = 5'h3 == _GEN_1115 ? 8'h0 : _GEN_1198; // @[CharOutput.scala 115:{23,23}]
  wire [7:0] _GEN_1200 = 5'h4 == _GEN_1115 ? 8'h6c : _GEN_1199; // @[CharOutput.scala 115:{23,23}]
  wire [7:0] _GEN_1201 = 5'h5 == _GEN_1115 ? 8'h0 : _GEN_1200; // @[CharOutput.scala 115:{23,23}]
  wire [7:0] _GEN_1202 = 5'h6 == _GEN_1115 ? 8'h0 : _GEN_1201; // @[CharOutput.scala 115:{23,23}]
  wire [7:0] _GEN_1203 = 5'h7 == _GEN_1115 ? 8'h0 : _GEN_1202; // @[CharOutput.scala 115:{23,23}]
  wire [7:0] _GEN_1204 = 5'h8 == _GEN_1115 ? 8'h72 : _GEN_1203; // @[CharOutput.scala 115:{23,23}]
  wire [7:0] _GEN_1205 = 5'h9 == _GEN_1115 ? 8'h0 : _GEN_1204; // @[CharOutput.scala 115:{23,23}]
  wire [7:0] _GEN_1206 = 5'ha == _GEN_1115 ? 8'h6e : _GEN_1205; // @[CharOutput.scala 115:{23,23}]
  wire [7:0] _GEN_1207 = 5'hb == _GEN_1115 ? 8'h0 : _GEN_1206; // @[CharOutput.scala 115:{23,23}]
  wire [7:0] _GEN_1208 = 5'hc == _GEN_1115 ? 8'h65 : _GEN_1207; // @[CharOutput.scala 115:{23,23}]
  wire [7:0] _GEN_1209 = 5'hd == _GEN_1115 ? 8'h72 : _GEN_1208; // @[CharOutput.scala 115:{23,23}]
  wire [7:0] _GEN_1210 = 5'he == _GEN_1115 ? 8'h6f : _GEN_1209; // @[CharOutput.scala 115:{23,23}]
  wire [7:0] _GEN_1211 = 5'hf == _GEN_1115 ? 8'h65 : _GEN_1210; // @[CharOutput.scala 115:{23,23}]
  wire [7:0] _GEN_1212 = 5'h10 == _GEN_1115 ? 8'h70 : _GEN_1211; // @[CharOutput.scala 115:{23,23}]
  wire [7:0] _GEN_1213 = 5'h11 == _GEN_1115 ? 8'h0 : _GEN_1212; // @[CharOutput.scala 115:{23,23}]
  wire [7:0] _GEN_1214 = 5'h12 == _GEN_1115 ? 8'h6e : _GEN_1213; // @[CharOutput.scala 115:{23,23}]
  wire [7:0] current_ascii_array_4 = 5'h13 == _GEN_1115 ? 8'h6e : _GEN_1214; // @[CharOutput.scala 115:{23,23}]
  wire [7:0] _GEN_1218 = 5'h2 == _GEN_1115 ? 8'h0 : 8'h6c; // @[CharOutput.scala 115:{23,23}]
  wire [7:0] _GEN_1219 = 5'h3 == _GEN_1115 ? 8'h0 : _GEN_1218; // @[CharOutput.scala 115:{23,23}]
  wire [7:0] _GEN_1220 = 5'h4 == _GEN_1115 ? 8'h65 : _GEN_1219; // @[CharOutput.scala 115:{23,23}]
  wire [7:0] _GEN_1221 = 5'h5 == _GEN_1115 ? 8'h0 : _GEN_1220; // @[CharOutput.scala 115:{23,23}]
  wire [7:0] _GEN_1222 = 5'h6 == _GEN_1115 ? 8'h0 : _GEN_1221; // @[CharOutput.scala 115:{23,23}]
  wire [7:0] _GEN_1223 = 5'h7 == _GEN_1115 ? 8'h0 : _GEN_1222; // @[CharOutput.scala 115:{23,23}]
  wire [7:0] _GEN_1224 = 5'h8 == _GEN_1115 ? 8'h0 : _GEN_1223; // @[CharOutput.scala 115:{23,23}]
  wire [7:0] _GEN_1225 = 5'h9 == _GEN_1115 ? 8'h0 : _GEN_1224; // @[CharOutput.scala 115:{23,23}]
  wire [7:0] _GEN_1226 = 5'ha == _GEN_1115 ? 8'h67 : _GEN_1225; // @[CharOutput.scala 115:{23,23}]
  wire [7:0] _GEN_1227 = 5'hb == _GEN_1115 ? 8'h0 : _GEN_1226; // @[CharOutput.scala 115:{23,23}]
  wire [7:0] _GEN_1228 = 5'hc == _GEN_1115 ? 8'h0 : _GEN_1227; // @[CharOutput.scala 115:{23,23}]
  wire [7:0] _GEN_1229 = 5'hd == _GEN_1115 ? 8'h62 : _GEN_1228; // @[CharOutput.scala 115:{23,23}]
  wire [7:0] _GEN_1230 = 5'he == _GEN_1115 ? 8'h6e : _GEN_1229; // @[CharOutput.scala 115:{23,23}]
  wire [7:0] _GEN_1231 = 5'hf == _GEN_1115 ? 8'h64 : _GEN_1230; // @[CharOutput.scala 115:{23,23}]
  wire [7:0] _GEN_1232 = 5'h10 == _GEN_1115 ? 8'h0 : _GEN_1231; // @[CharOutput.scala 115:{23,23}]
  wire [7:0] _GEN_1233 = 5'h11 == _GEN_1115 ? 8'h0 : _GEN_1232; // @[CharOutput.scala 115:{23,23}]
  wire [7:0] _GEN_1234 = 5'h12 == _GEN_1115 ? 8'h0 : _GEN_1233; // @[CharOutput.scala 115:{23,23}]
  wire [7:0] current_ascii_array_5 = 5'h13 == _GEN_1115 ? 8'h69 : _GEN_1234; // @[CharOutput.scala 115:{23,23}]
  wire [7:0] _GEN_1237 = 5'h1 == _GEN_1115 ? 8'h65 : 8'h61; // @[CharOutput.scala 115:{23,23}]
  wire [7:0] _GEN_1238 = 5'h2 == _GEN_1115 ? 8'h0 : _GEN_1237; // @[CharOutput.scala 115:{23,23}]
  wire [7:0] _GEN_1239 = 5'h3 == _GEN_1115 ? 8'h0 : _GEN_1238; // @[CharOutput.scala 115:{23,23}]
  wire [7:0] _GEN_1240 = 5'h4 == _GEN_1115 ? 8'h0 : _GEN_1239; // @[CharOutput.scala 115:{23,23}]
  wire [7:0] _GEN_1241 = 5'h5 == _GEN_1115 ? 8'h0 : _GEN_1240; // @[CharOutput.scala 115:{23,23}]
  wire [7:0] _GEN_1242 = 5'h6 == _GEN_1115 ? 8'h0 : _GEN_1241; // @[CharOutput.scala 115:{23,23}]
  wire [7:0] _GEN_1243 = 5'h7 == _GEN_1115 ? 8'h0 : _GEN_1242; // @[CharOutput.scala 115:{23,23}]
  wire [7:0] _GEN_1244 = 5'h8 == _GEN_1115 ? 8'h0 : _GEN_1243; // @[CharOutput.scala 115:{23,23}]
  wire [7:0] _GEN_1245 = 5'h9 == _GEN_1115 ? 8'h0 : _GEN_1244; // @[CharOutput.scala 115:{23,23}]
  wire [7:0] _GEN_1246 = 5'ha == _GEN_1115 ? 8'h74 : _GEN_1245; // @[CharOutput.scala 115:{23,23}]
  wire [7:0] _GEN_1247 = 5'hb == _GEN_1115 ? 8'h0 : _GEN_1246; // @[CharOutput.scala 115:{23,23}]
  wire [7:0] _GEN_1248 = 5'hc == _GEN_1115 ? 8'h0 : _GEN_1247; // @[CharOutput.scala 115:{23,23}]
  wire [7:0] _GEN_1249 = 5'hd == _GEN_1115 ? 8'h69 : _GEN_1248; // @[CharOutput.scala 115:{23,23}]
  wire [7:0] _GEN_1250 = 5'he == _GEN_1115 ? 8'h0 : _GEN_1249; // @[CharOutput.scala 115:{23,23}]
  wire [7:0] _GEN_1251 = 5'hf == _GEN_1115 ? 8'h70 : _GEN_1250; // @[CharOutput.scala 115:{23,23}]
  wire [7:0] _GEN_1252 = 5'h10 == _GEN_1115 ? 8'h0 : _GEN_1251; // @[CharOutput.scala 115:{23,23}]
  wire [7:0] _GEN_1253 = 5'h11 == _GEN_1115 ? 8'h0 : _GEN_1252; // @[CharOutput.scala 115:{23,23}]
  wire [7:0] _GEN_1254 = 5'h12 == _GEN_1115 ? 8'h0 : _GEN_1253; // @[CharOutput.scala 115:{23,23}]
  wire [7:0] current_ascii_array_6 = 5'h13 == _GEN_1115 ? 8'h74 : _GEN_1254; // @[CharOutput.scala 115:{23,23}]
  wire [7:0] _GEN_1257 = 5'h1 == _GEN_1115 ? 8'h0 : 8'h6e; // @[CharOutput.scala 115:{23,23}]
  wire [7:0] _GEN_1258 = 5'h2 == _GEN_1115 ? 8'h0 : _GEN_1257; // @[CharOutput.scala 115:{23,23}]
  wire [7:0] _GEN_1259 = 5'h3 == _GEN_1115 ? 8'h0 : _GEN_1258; // @[CharOutput.scala 115:{23,23}]
  wire [7:0] _GEN_1260 = 5'h4 == _GEN_1115 ? 8'h0 : _GEN_1259; // @[CharOutput.scala 115:{23,23}]
  wire [7:0] _GEN_1261 = 5'h5 == _GEN_1115 ? 8'h0 : _GEN_1260; // @[CharOutput.scala 115:{23,23}]
  wire [7:0] _GEN_1262 = 5'h6 == _GEN_1115 ? 8'h0 : _GEN_1261; // @[CharOutput.scala 115:{23,23}]
  wire [7:0] _GEN_1263 = 5'h7 == _GEN_1115 ? 8'h0 : _GEN_1262; // @[CharOutput.scala 115:{23,23}]
  wire [7:0] _GEN_1264 = 5'h8 == _GEN_1115 ? 8'h0 : _GEN_1263; // @[CharOutput.scala 115:{23,23}]
  wire [7:0] _GEN_1265 = 5'h9 == _GEN_1115 ? 8'h0 : _GEN_1264; // @[CharOutput.scala 115:{23,23}]
  wire [7:0] _GEN_1266 = 5'ha == _GEN_1115 ? 8'h61 : _GEN_1265; // @[CharOutput.scala 115:{23,23}]
  wire [7:0] _GEN_1267 = 5'hb == _GEN_1115 ? 8'h0 : _GEN_1266; // @[CharOutput.scala 115:{23,23}]
  wire [7:0] _GEN_1268 = 5'hc == _GEN_1115 ? 8'h0 : _GEN_1267; // @[CharOutput.scala 115:{23,23}]
  wire [7:0] _GEN_1269 = 5'hd == _GEN_1115 ? 8'h6b : _GEN_1268; // @[CharOutput.scala 115:{23,23}]
  wire [7:0] _GEN_1270 = 5'he == _GEN_1115 ? 8'h0 : _GEN_1269; // @[CharOutput.scala 115:{23,23}]
  wire [7:0] _GEN_1271 = 5'hf == _GEN_1115 ? 8'h6c : _GEN_1270; // @[CharOutput.scala 115:{23,23}]
  wire [7:0] _GEN_1272 = 5'h10 == _GEN_1115 ? 8'h0 : _GEN_1271; // @[CharOutput.scala 115:{23,23}]
  wire [7:0] _GEN_1273 = 5'h11 == _GEN_1115 ? 8'h0 : _GEN_1272; // @[CharOutput.scala 115:{23,23}]
  wire [7:0] _GEN_1274 = 5'h12 == _GEN_1115 ? 8'h0 : _GEN_1273; // @[CharOutput.scala 115:{23,23}]
  wire [7:0] current_ascii_array_7 = 5'h13 == _GEN_1115 ? 8'h6f : _GEN_1274; // @[CharOutput.scala 115:{23,23}]
  wire [7:0] _GEN_1277 = 5'h1 == _GEN_1115 ? 8'h0 : 8'h65; // @[CharOutput.scala 115:{23,23}]
  wire [7:0] _GEN_1278 = 5'h2 == _GEN_1115 ? 8'h0 : _GEN_1277; // @[CharOutput.scala 115:{23,23}]
  wire [7:0] _GEN_1279 = 5'h3 == _GEN_1115 ? 8'h0 : _GEN_1278; // @[CharOutput.scala 115:{23,23}]
  wire [7:0] _GEN_1280 = 5'h4 == _GEN_1115 ? 8'h0 : _GEN_1279; // @[CharOutput.scala 115:{23,23}]
  wire [7:0] _GEN_1281 = 5'h5 == _GEN_1115 ? 8'h0 : _GEN_1280; // @[CharOutput.scala 115:{23,23}]
  wire [7:0] _GEN_1282 = 5'h6 == _GEN_1115 ? 8'h0 : _GEN_1281; // @[CharOutput.scala 115:{23,23}]
  wire [7:0] _GEN_1283 = 5'h7 == _GEN_1115 ? 8'h0 : _GEN_1282; // @[CharOutput.scala 115:{23,23}]
  wire [7:0] _GEN_1284 = 5'h8 == _GEN_1115 ? 8'h0 : _GEN_1283; // @[CharOutput.scala 115:{23,23}]
  wire [7:0] _GEN_1285 = 5'h9 == _GEN_1115 ? 8'h0 : _GEN_1284; // @[CharOutput.scala 115:{23,23}]
  wire [7:0] _GEN_1286 = 5'ha == _GEN_1115 ? 8'h62 : _GEN_1285; // @[CharOutput.scala 115:{23,23}]
  wire [7:0] _GEN_1287 = 5'hb == _GEN_1115 ? 8'h0 : _GEN_1286; // @[CharOutput.scala 115:{23,23}]
  wire [7:0] _GEN_1288 = 5'hc == _GEN_1115 ? 8'h0 : _GEN_1287; // @[CharOutput.scala 115:{23,23}]
  wire [7:0] _GEN_1289 = 5'hd == _GEN_1115 ? 8'h65 : _GEN_1288; // @[CharOutput.scala 115:{23,23}]
  wire [7:0] _GEN_1290 = 5'he == _GEN_1115 ? 8'h0 : _GEN_1289; // @[CharOutput.scala 115:{23,23}]
  wire [7:0] _GEN_1291 = 5'hf == _GEN_1115 ? 8'h61 : _GEN_1290; // @[CharOutput.scala 115:{23,23}]
  wire [7:0] _GEN_1292 = 5'h10 == _GEN_1115 ? 8'h0 : _GEN_1291; // @[CharOutput.scala 115:{23,23}]
  wire [7:0] _GEN_1293 = 5'h11 == _GEN_1115 ? 8'h0 : _GEN_1292; // @[CharOutput.scala 115:{23,23}]
  wire [7:0] _GEN_1294 = 5'h12 == _GEN_1115 ? 8'h0 : _GEN_1293; // @[CharOutput.scala 115:{23,23}]
  wire [7:0] current_ascii_array_8 = 5'h13 == _GEN_1115 ? 8'h72 : _GEN_1294; // @[CharOutput.scala 115:{23,23}]
  wire [7:0] _GEN_1306 = 5'ha == _GEN_1115 ? 8'h6c : 8'h0; // @[CharOutput.scala 115:{23,23}]
  wire [7:0] _GEN_1307 = 5'hb == _GEN_1115 ? 8'h0 : _GEN_1306; // @[CharOutput.scala 115:{23,23}]
  wire [7:0] _GEN_1308 = 5'hc == _GEN_1115 ? 8'h0 : _GEN_1307; // @[CharOutput.scala 115:{23,23}]
  wire [7:0] _GEN_1309 = 5'hd == _GEN_1115 ? 8'h0 : _GEN_1308; // @[CharOutput.scala 115:{23,23}]
  wire [7:0] _GEN_1310 = 5'he == _GEN_1115 ? 8'h0 : _GEN_1309; // @[CharOutput.scala 115:{23,23}]
  wire [7:0] _GEN_1311 = 5'hf == _GEN_1115 ? 8'h6e : _GEN_1310; // @[CharOutput.scala 115:{23,23}]
  wire [7:0] _GEN_1312 = 5'h10 == _GEN_1115 ? 8'h0 : _GEN_1311; // @[CharOutput.scala 115:{23,23}]
  wire [7:0] _GEN_1313 = 5'h11 == _GEN_1115 ? 8'h0 : _GEN_1312; // @[CharOutput.scala 115:{23,23}]
  wire [7:0] _GEN_1314 = 5'h12 == _GEN_1115 ? 8'h0 : _GEN_1313; // @[CharOutput.scala 115:{23,23}]
  wire [7:0] current_ascii_array_9 = 5'h13 == _GEN_1115 ? 8'h0 : _GEN_1314; // @[CharOutput.scala 115:{23,23}]
  wire [7:0] _GEN_1326 = 5'ha == _GEN_1115 ? 8'h65 : 8'h0; // @[CharOutput.scala 115:{23,23}]
  wire [7:0] _GEN_1327 = 5'hb == _GEN_1115 ? 8'h0 : _GEN_1326; // @[CharOutput.scala 115:{23,23}]
  wire [7:0] _GEN_1328 = 5'hc == _GEN_1115 ? 8'h0 : _GEN_1327; // @[CharOutput.scala 115:{23,23}]
  wire [7:0] _GEN_1329 = 5'hd == _GEN_1115 ? 8'h0 : _GEN_1328; // @[CharOutput.scala 115:{23,23}]
  wire [7:0] _GEN_1330 = 5'he == _GEN_1115 ? 8'h0 : _GEN_1329; // @[CharOutput.scala 115:{23,23}]
  wire [7:0] _GEN_1331 = 5'hf == _GEN_1115 ? 8'h74 : _GEN_1330; // @[CharOutput.scala 115:{23,23}]
  wire [7:0] _GEN_1332 = 5'h10 == _GEN_1115 ? 8'h0 : _GEN_1331; // @[CharOutput.scala 115:{23,23}]
  wire [7:0] _GEN_1333 = 5'h11 == _GEN_1115 ? 8'h0 : _GEN_1332; // @[CharOutput.scala 115:{23,23}]
  wire [7:0] _GEN_1334 = 5'h12 == _GEN_1115 ? 8'h0 : _GEN_1333; // @[CharOutput.scala 115:{23,23}]
  wire [7:0] current_ascii_array_10 = 5'h13 == _GEN_1115 ? 8'h0 : _GEN_1334; // @[CharOutput.scala 115:{23,23}]
  wire [3:0] _GEN_1337 = 3'h1 == obj_choose ? char_index_1 : char_index_0; // @[CharOutput.scala 116:{17,17}]
  wire [3:0] _GEN_1338 = 3'h2 == obj_choose ? char_index_2 : _GEN_1337; // @[CharOutput.scala 116:{17,17}]
  wire [3:0] _GEN_1339 = 3'h3 == obj_choose ? char_index_3 : _GEN_1338; // @[CharOutput.scala 116:{17,17}]
  wire [3:0] _GEN_1340 = 3'h4 == obj_choose ? char_index_4 : _GEN_1339; // @[CharOutput.scala 116:{17,17}]
  wire [7:0] _GEN_1342 = 4'h1 == _GEN_1340 ? current_ascii_array_1 : current_ascii_array_0; // @[CharOutput.scala 116:{17,17}]
  wire [7:0] _GEN_1343 = 4'h2 == _GEN_1340 ? current_ascii_array_2 : _GEN_1342; // @[CharOutput.scala 116:{17,17}]
  wire [7:0] _GEN_1344 = 4'h3 == _GEN_1340 ? current_ascii_array_3 : _GEN_1343; // @[CharOutput.scala 116:{17,17}]
  wire [7:0] _GEN_1345 = 4'h4 == _GEN_1340 ? current_ascii_array_4 : _GEN_1344; // @[CharOutput.scala 116:{17,17}]
  wire [7:0] _GEN_1346 = 4'h5 == _GEN_1340 ? current_ascii_array_5 : _GEN_1345; // @[CharOutput.scala 116:{17,17}]
  wire [7:0] _GEN_1347 = 4'h6 == _GEN_1340 ? current_ascii_array_6 : _GEN_1346; // @[CharOutput.scala 116:{17,17}]
  wire [7:0] _GEN_1348 = 4'h7 == _GEN_1340 ? current_ascii_array_7 : _GEN_1347; // @[CharOutput.scala 116:{17,17}]
  wire [7:0] _GEN_1349 = 4'h8 == _GEN_1340 ? current_ascii_array_8 : _GEN_1348; // @[CharOutput.scala 116:{17,17}]
  wire [7:0] _GEN_1350 = 4'h9 == _GEN_1340 ? current_ascii_array_9 : _GEN_1349; // @[CharOutput.scala 116:{17,17}]
  wire [7:0] current_ascii = 4'ha == _GEN_1340 ? current_ascii_array_10 : _GEN_1350; // @[CharOutput.scala 116:{17,17}]
  wire [12:0] char_baseaddr_lut_0 = {{7'd0}, _char_baseaddr_lut_T}; // @[CharOutput.scala 110:{34,34}]
  wire [12:0] char_baseaddr_lut_1 = {{7'd0}, _char_baseaddr_lut_T_1}; // @[CharOutput.scala 110:{34,34}]
  wire [12:0] _GEN_1353 = 8'h1 == current_ascii ? char_baseaddr_lut_1 : char_baseaddr_lut_0; // @[CharOutput.scala 118:{17,17}]
  wire [12:0] char_baseaddr_lut_2 = {{6'd0}, _char_baseaddr_lut_T_2}; // @[CharOutput.scala 110:{34,34}]
  wire [12:0] _GEN_1354 = 8'h2 == current_ascii ? char_baseaddr_lut_2 : _GEN_1353; // @[CharOutput.scala 118:{17,17}]
  wire [12:0] char_baseaddr_lut_3 = {{6'd0}, _char_baseaddr_lut_T_3}; // @[CharOutput.scala 110:{34,34}]
  wire [12:0] _GEN_1355 = 8'h3 == current_ascii ? char_baseaddr_lut_3 : _GEN_1354; // @[CharOutput.scala 118:{17,17}]
  wire [12:0] char_baseaddr_lut_4 = {{5'd0}, _char_baseaddr_lut_T_4}; // @[CharOutput.scala 110:{34,34}]
  wire [12:0] _GEN_1356 = 8'h4 == current_ascii ? char_baseaddr_lut_4 : _GEN_1355; // @[CharOutput.scala 118:{17,17}]
  wire [12:0] char_baseaddr_lut_5 = {{5'd0}, _char_baseaddr_lut_T_5}; // @[CharOutput.scala 110:{34,34}]
  wire [12:0] _GEN_1357 = 8'h5 == current_ascii ? char_baseaddr_lut_5 : _GEN_1356; // @[CharOutput.scala 118:{17,17}]
  wire [12:0] char_baseaddr_lut_6 = {{5'd0}, _char_baseaddr_lut_T_6}; // @[CharOutput.scala 110:{34,34}]
  wire [12:0] _GEN_1358 = 8'h6 == current_ascii ? char_baseaddr_lut_6 : _GEN_1357; // @[CharOutput.scala 118:{17,17}]
  wire [12:0] char_baseaddr_lut_7 = {{5'd0}, _char_baseaddr_lut_T_7}; // @[CharOutput.scala 110:{34,34}]
  wire [12:0] _GEN_1359 = 8'h7 == current_ascii ? char_baseaddr_lut_7 : _GEN_1358; // @[CharOutput.scala 118:{17,17}]
  wire [12:0] char_baseaddr_lut_8 = {{4'd0}, _char_baseaddr_lut_T_8}; // @[CharOutput.scala 110:{34,34}]
  wire [12:0] _GEN_1360 = 8'h8 == current_ascii ? char_baseaddr_lut_8 : _GEN_1359; // @[CharOutput.scala 118:{17,17}]
  wire [12:0] char_baseaddr_lut_9 = {{4'd0}, _char_baseaddr_lut_T_9}; // @[CharOutput.scala 110:{34,34}]
  wire [12:0] _GEN_1361 = 8'h9 == current_ascii ? char_baseaddr_lut_9 : _GEN_1360; // @[CharOutput.scala 118:{17,17}]
  wire [12:0] char_baseaddr_lut_10 = {{4'd0}, _char_baseaddr_lut_T_10}; // @[CharOutput.scala 110:{34,34}]
  wire [12:0] _GEN_1362 = 8'ha == current_ascii ? char_baseaddr_lut_10 : _GEN_1361; // @[CharOutput.scala 118:{17,17}]
  wire [12:0] char_baseaddr_lut_11 = {{4'd0}, _char_baseaddr_lut_T_11}; // @[CharOutput.scala 110:{34,34}]
  wire [12:0] _GEN_1363 = 8'hb == current_ascii ? char_baseaddr_lut_11 : _GEN_1362; // @[CharOutput.scala 118:{17,17}]
  wire [12:0] char_baseaddr_lut_12 = {{4'd0}, _char_baseaddr_lut_T_12}; // @[CharOutput.scala 110:{34,34}]
  wire [12:0] _GEN_1364 = 8'hc == current_ascii ? char_baseaddr_lut_12 : _GEN_1363; // @[CharOutput.scala 118:{17,17}]
  wire [12:0] char_baseaddr_lut_13 = {{4'd0}, _char_baseaddr_lut_T_13}; // @[CharOutput.scala 110:{34,34}]
  wire [12:0] _GEN_1365 = 8'hd == current_ascii ? char_baseaddr_lut_13 : _GEN_1364; // @[CharOutput.scala 118:{17,17}]
  wire [12:0] char_baseaddr_lut_14 = {{4'd0}, _char_baseaddr_lut_T_14}; // @[CharOutput.scala 110:{34,34}]
  wire [12:0] _GEN_1366 = 8'he == current_ascii ? char_baseaddr_lut_14 : _GEN_1365; // @[CharOutput.scala 118:{17,17}]
  wire [12:0] char_baseaddr_lut_15 = {{4'd0}, _char_baseaddr_lut_T_15}; // @[CharOutput.scala 110:{34,34}]
  wire [12:0] _GEN_1367 = 8'hf == current_ascii ? char_baseaddr_lut_15 : _GEN_1366; // @[CharOutput.scala 118:{17,17}]
  wire [12:0] char_baseaddr_lut_16 = {{3'd0}, _char_baseaddr_lut_T_16}; // @[CharOutput.scala 110:{34,34}]
  wire [12:0] _GEN_1368 = 8'h10 == current_ascii ? char_baseaddr_lut_16 : _GEN_1367; // @[CharOutput.scala 118:{17,17}]
  wire [12:0] char_baseaddr_lut_17 = {{3'd0}, _char_baseaddr_lut_T_17}; // @[CharOutput.scala 110:{34,34}]
  wire [12:0] _GEN_1369 = 8'h11 == current_ascii ? char_baseaddr_lut_17 : _GEN_1368; // @[CharOutput.scala 118:{17,17}]
  wire [12:0] char_baseaddr_lut_18 = {{3'd0}, _char_baseaddr_lut_T_18}; // @[CharOutput.scala 110:{34,34}]
  wire [12:0] _GEN_1370 = 8'h12 == current_ascii ? char_baseaddr_lut_18 : _GEN_1369; // @[CharOutput.scala 118:{17,17}]
  wire [12:0] char_baseaddr_lut_19 = {{3'd0}, _char_baseaddr_lut_T_19}; // @[CharOutput.scala 110:{34,34}]
  wire [12:0] _GEN_1371 = 8'h13 == current_ascii ? char_baseaddr_lut_19 : _GEN_1370; // @[CharOutput.scala 118:{17,17}]
  wire [12:0] char_baseaddr_lut_20 = {{3'd0}, _char_baseaddr_lut_T_20}; // @[CharOutput.scala 110:{34,34}]
  wire [12:0] _GEN_1372 = 8'h14 == current_ascii ? char_baseaddr_lut_20 : _GEN_1371; // @[CharOutput.scala 118:{17,17}]
  wire [12:0] char_baseaddr_lut_21 = {{3'd0}, _char_baseaddr_lut_T_21}; // @[CharOutput.scala 110:{34,34}]
  wire [12:0] _GEN_1373 = 8'h15 == current_ascii ? char_baseaddr_lut_21 : _GEN_1372; // @[CharOutput.scala 118:{17,17}]
  wire [12:0] char_baseaddr_lut_22 = {{3'd0}, _char_baseaddr_lut_T_22}; // @[CharOutput.scala 110:{34,34}]
  wire [12:0] _GEN_1374 = 8'h16 == current_ascii ? char_baseaddr_lut_22 : _GEN_1373; // @[CharOutput.scala 118:{17,17}]
  wire [12:0] char_baseaddr_lut_23 = {{3'd0}, _char_baseaddr_lut_T_23}; // @[CharOutput.scala 110:{34,34}]
  wire [12:0] _GEN_1375 = 8'h17 == current_ascii ? char_baseaddr_lut_23 : _GEN_1374; // @[CharOutput.scala 118:{17,17}]
  wire [12:0] char_baseaddr_lut_24 = {{3'd0}, _char_baseaddr_lut_T_24}; // @[CharOutput.scala 110:{34,34}]
  wire [12:0] _GEN_1376 = 8'h18 == current_ascii ? char_baseaddr_lut_24 : _GEN_1375; // @[CharOutput.scala 118:{17,17}]
  wire [12:0] char_baseaddr_lut_25 = {{3'd0}, _char_baseaddr_lut_T_25}; // @[CharOutput.scala 110:{34,34}]
  wire [12:0] _GEN_1377 = 8'h19 == current_ascii ? char_baseaddr_lut_25 : _GEN_1376; // @[CharOutput.scala 118:{17,17}]
  wire [12:0] char_baseaddr_lut_26 = {{3'd0}, _char_baseaddr_lut_T_26}; // @[CharOutput.scala 110:{34,34}]
  wire [12:0] _GEN_1378 = 8'h1a == current_ascii ? char_baseaddr_lut_26 : _GEN_1377; // @[CharOutput.scala 118:{17,17}]
  wire [12:0] char_baseaddr_lut_27 = {{3'd0}, _char_baseaddr_lut_T_27}; // @[CharOutput.scala 110:{34,34}]
  wire [12:0] _GEN_1379 = 8'h1b == current_ascii ? char_baseaddr_lut_27 : _GEN_1378; // @[CharOutput.scala 118:{17,17}]
  wire [12:0] char_baseaddr_lut_28 = {{3'd0}, _char_baseaddr_lut_T_28}; // @[CharOutput.scala 110:{34,34}]
  wire [12:0] _GEN_1380 = 8'h1c == current_ascii ? char_baseaddr_lut_28 : _GEN_1379; // @[CharOutput.scala 118:{17,17}]
  wire [12:0] char_baseaddr_lut_29 = {{3'd0}, _char_baseaddr_lut_T_29}; // @[CharOutput.scala 110:{34,34}]
  wire [12:0] _GEN_1381 = 8'h1d == current_ascii ? char_baseaddr_lut_29 : _GEN_1380; // @[CharOutput.scala 118:{17,17}]
  wire [12:0] char_baseaddr_lut_30 = {{3'd0}, _char_baseaddr_lut_T_30}; // @[CharOutput.scala 110:{34,34}]
  wire [12:0] _GEN_1382 = 8'h1e == current_ascii ? char_baseaddr_lut_30 : _GEN_1381; // @[CharOutput.scala 118:{17,17}]
  wire [12:0] char_baseaddr_lut_31 = {{3'd0}, _char_baseaddr_lut_T_31}; // @[CharOutput.scala 110:{34,34}]
  wire [12:0] _GEN_1383 = 8'h1f == current_ascii ? char_baseaddr_lut_31 : _GEN_1382; // @[CharOutput.scala 118:{17,17}]
  wire [12:0] char_baseaddr_lut_32 = {{2'd0}, _char_baseaddr_lut_T_32}; // @[CharOutput.scala 110:{34,34}]
  wire [12:0] _GEN_1384 = 8'h20 == current_ascii ? char_baseaddr_lut_32 : _GEN_1383; // @[CharOutput.scala 118:{17,17}]
  wire [12:0] char_baseaddr_lut_33 = {{2'd0}, _char_baseaddr_lut_T_33}; // @[CharOutput.scala 110:{34,34}]
  wire [12:0] _GEN_1385 = 8'h21 == current_ascii ? char_baseaddr_lut_33 : _GEN_1384; // @[CharOutput.scala 118:{17,17}]
  wire [12:0] char_baseaddr_lut_34 = {{2'd0}, _char_baseaddr_lut_T_34}; // @[CharOutput.scala 110:{34,34}]
  wire [12:0] _GEN_1386 = 8'h22 == current_ascii ? char_baseaddr_lut_34 : _GEN_1385; // @[CharOutput.scala 118:{17,17}]
  wire [12:0] char_baseaddr_lut_35 = {{2'd0}, _char_baseaddr_lut_T_35}; // @[CharOutput.scala 110:{34,34}]
  wire [12:0] _GEN_1387 = 8'h23 == current_ascii ? char_baseaddr_lut_35 : _GEN_1386; // @[CharOutput.scala 118:{17,17}]
  wire [12:0] char_baseaddr_lut_36 = {{2'd0}, _char_baseaddr_lut_T_36}; // @[CharOutput.scala 110:{34,34}]
  wire [12:0] _GEN_1388 = 8'h24 == current_ascii ? char_baseaddr_lut_36 : _GEN_1387; // @[CharOutput.scala 118:{17,17}]
  wire [12:0] char_baseaddr_lut_37 = {{2'd0}, _char_baseaddr_lut_T_37}; // @[CharOutput.scala 110:{34,34}]
  wire [12:0] _GEN_1389 = 8'h25 == current_ascii ? char_baseaddr_lut_37 : _GEN_1388; // @[CharOutput.scala 118:{17,17}]
  wire [12:0] char_baseaddr_lut_38 = {{2'd0}, _char_baseaddr_lut_T_38}; // @[CharOutput.scala 110:{34,34}]
  wire [12:0] _GEN_1390 = 8'h26 == current_ascii ? char_baseaddr_lut_38 : _GEN_1389; // @[CharOutput.scala 118:{17,17}]
  wire [12:0] char_baseaddr_lut_39 = {{2'd0}, _char_baseaddr_lut_T_39}; // @[CharOutput.scala 110:{34,34}]
  wire [12:0] _GEN_1391 = 8'h27 == current_ascii ? char_baseaddr_lut_39 : _GEN_1390; // @[CharOutput.scala 118:{17,17}]
  wire [12:0] char_baseaddr_lut_40 = {{2'd0}, _char_baseaddr_lut_T_40}; // @[CharOutput.scala 110:{34,34}]
  wire [12:0] _GEN_1392 = 8'h28 == current_ascii ? char_baseaddr_lut_40 : _GEN_1391; // @[CharOutput.scala 118:{17,17}]
  wire [12:0] char_baseaddr_lut_41 = {{2'd0}, _char_baseaddr_lut_T_41}; // @[CharOutput.scala 110:{34,34}]
  wire [12:0] _GEN_1393 = 8'h29 == current_ascii ? char_baseaddr_lut_41 : _GEN_1392; // @[CharOutput.scala 118:{17,17}]
  wire [12:0] char_baseaddr_lut_42 = {{2'd0}, _char_baseaddr_lut_T_42}; // @[CharOutput.scala 110:{34,34}]
  wire [12:0] _GEN_1394 = 8'h2a == current_ascii ? char_baseaddr_lut_42 : _GEN_1393; // @[CharOutput.scala 118:{17,17}]
  wire [12:0] char_baseaddr_lut_43 = {{2'd0}, _char_baseaddr_lut_T_43}; // @[CharOutput.scala 110:{34,34}]
  wire [12:0] _GEN_1395 = 8'h2b == current_ascii ? char_baseaddr_lut_43 : _GEN_1394; // @[CharOutput.scala 118:{17,17}]
  wire [12:0] char_baseaddr_lut_44 = {{2'd0}, _char_baseaddr_lut_T_44}; // @[CharOutput.scala 110:{34,34}]
  wire [12:0] _GEN_1396 = 8'h2c == current_ascii ? char_baseaddr_lut_44 : _GEN_1395; // @[CharOutput.scala 118:{17,17}]
  wire [12:0] char_baseaddr_lut_45 = {{2'd0}, _char_baseaddr_lut_T_45}; // @[CharOutput.scala 110:{34,34}]
  wire [12:0] _GEN_1397 = 8'h2d == current_ascii ? char_baseaddr_lut_45 : _GEN_1396; // @[CharOutput.scala 118:{17,17}]
  wire [12:0] char_baseaddr_lut_46 = {{2'd0}, _char_baseaddr_lut_T_46}; // @[CharOutput.scala 110:{34,34}]
  wire [12:0] _GEN_1398 = 8'h2e == current_ascii ? char_baseaddr_lut_46 : _GEN_1397; // @[CharOutput.scala 118:{17,17}]
  wire [12:0] char_baseaddr_lut_47 = {{2'd0}, _char_baseaddr_lut_T_47}; // @[CharOutput.scala 110:{34,34}]
  wire [12:0] _GEN_1399 = 8'h2f == current_ascii ? char_baseaddr_lut_47 : _GEN_1398; // @[CharOutput.scala 118:{17,17}]
  wire [12:0] char_baseaddr_lut_48 = {{2'd0}, _char_baseaddr_lut_T_48}; // @[CharOutput.scala 110:{34,34}]
  wire [12:0] _GEN_1400 = 8'h30 == current_ascii ? char_baseaddr_lut_48 : _GEN_1399; // @[CharOutput.scala 118:{17,17}]
  wire [12:0] char_baseaddr_lut_49 = {{2'd0}, _char_baseaddr_lut_T_49}; // @[CharOutput.scala 110:{34,34}]
  wire [12:0] _GEN_1401 = 8'h31 == current_ascii ? char_baseaddr_lut_49 : _GEN_1400; // @[CharOutput.scala 118:{17,17}]
  wire [12:0] char_baseaddr_lut_50 = {{2'd0}, _char_baseaddr_lut_T_50}; // @[CharOutput.scala 110:{34,34}]
  wire [12:0] _GEN_1402 = 8'h32 == current_ascii ? char_baseaddr_lut_50 : _GEN_1401; // @[CharOutput.scala 118:{17,17}]
  wire [12:0] char_baseaddr_lut_51 = {{2'd0}, _char_baseaddr_lut_T_51}; // @[CharOutput.scala 110:{34,34}]
  wire [12:0] _GEN_1403 = 8'h33 == current_ascii ? char_baseaddr_lut_51 : _GEN_1402; // @[CharOutput.scala 118:{17,17}]
  wire [12:0] char_baseaddr_lut_52 = {{2'd0}, _char_baseaddr_lut_T_52}; // @[CharOutput.scala 110:{34,34}]
  wire [12:0] _GEN_1404 = 8'h34 == current_ascii ? char_baseaddr_lut_52 : _GEN_1403; // @[CharOutput.scala 118:{17,17}]
  wire [12:0] char_baseaddr_lut_53 = {{2'd0}, _char_baseaddr_lut_T_53}; // @[CharOutput.scala 110:{34,34}]
  wire [12:0] _GEN_1405 = 8'h35 == current_ascii ? char_baseaddr_lut_53 : _GEN_1404; // @[CharOutput.scala 118:{17,17}]
  wire [12:0] char_baseaddr_lut_54 = {{2'd0}, _char_baseaddr_lut_T_54}; // @[CharOutput.scala 110:{34,34}]
  wire [12:0] _GEN_1406 = 8'h36 == current_ascii ? char_baseaddr_lut_54 : _GEN_1405; // @[CharOutput.scala 118:{17,17}]
  wire [12:0] char_baseaddr_lut_55 = {{2'd0}, _char_baseaddr_lut_T_55}; // @[CharOutput.scala 110:{34,34}]
  wire [12:0] _GEN_1407 = 8'h37 == current_ascii ? char_baseaddr_lut_55 : _GEN_1406; // @[CharOutput.scala 118:{17,17}]
  wire [12:0] char_baseaddr_lut_56 = {{2'd0}, _char_baseaddr_lut_T_56}; // @[CharOutput.scala 110:{34,34}]
  wire [12:0] _GEN_1408 = 8'h38 == current_ascii ? char_baseaddr_lut_56 : _GEN_1407; // @[CharOutput.scala 118:{17,17}]
  wire [12:0] char_baseaddr_lut_57 = {{2'd0}, _char_baseaddr_lut_T_57}; // @[CharOutput.scala 110:{34,34}]
  wire [12:0] _GEN_1409 = 8'h39 == current_ascii ? char_baseaddr_lut_57 : _GEN_1408; // @[CharOutput.scala 118:{17,17}]
  wire [12:0] char_baseaddr_lut_58 = {{2'd0}, _char_baseaddr_lut_T_58}; // @[CharOutput.scala 110:{34,34}]
  wire [12:0] _GEN_1410 = 8'h3a == current_ascii ? char_baseaddr_lut_58 : _GEN_1409; // @[CharOutput.scala 118:{17,17}]
  wire [12:0] char_baseaddr_lut_59 = {{2'd0}, _char_baseaddr_lut_T_59}; // @[CharOutput.scala 110:{34,34}]
  wire [12:0] _GEN_1411 = 8'h3b == current_ascii ? char_baseaddr_lut_59 : _GEN_1410; // @[CharOutput.scala 118:{17,17}]
  wire [12:0] char_baseaddr_lut_60 = {{2'd0}, _char_baseaddr_lut_T_60}; // @[CharOutput.scala 110:{34,34}]
  wire [12:0] _GEN_1412 = 8'h3c == current_ascii ? char_baseaddr_lut_60 : _GEN_1411; // @[CharOutput.scala 118:{17,17}]
  wire [12:0] char_baseaddr_lut_61 = {{2'd0}, _char_baseaddr_lut_T_61}; // @[CharOutput.scala 110:{34,34}]
  wire [12:0] _GEN_1413 = 8'h3d == current_ascii ? char_baseaddr_lut_61 : _GEN_1412; // @[CharOutput.scala 118:{17,17}]
  wire [12:0] char_baseaddr_lut_62 = {{2'd0}, _char_baseaddr_lut_T_62}; // @[CharOutput.scala 110:{34,34}]
  wire [12:0] _GEN_1414 = 8'h3e == current_ascii ? char_baseaddr_lut_62 : _GEN_1413; // @[CharOutput.scala 118:{17,17}]
  wire [12:0] char_baseaddr_lut_63 = {{2'd0}, _char_baseaddr_lut_T_63}; // @[CharOutput.scala 110:{34,34}]
  wire [12:0] _GEN_1415 = 8'h3f == current_ascii ? char_baseaddr_lut_63 : _GEN_1414; // @[CharOutput.scala 118:{17,17}]
  wire [12:0] char_baseaddr_lut_64 = {{1'd0}, _char_baseaddr_lut_T_64}; // @[CharOutput.scala 110:{34,34}]
  wire [12:0] _GEN_1416 = 8'h40 == current_ascii ? char_baseaddr_lut_64 : _GEN_1415; // @[CharOutput.scala 118:{17,17}]
  wire [12:0] char_baseaddr_lut_65 = {{1'd0}, _char_baseaddr_lut_T_65}; // @[CharOutput.scala 110:{34,34}]
  wire [12:0] _GEN_1417 = 8'h41 == current_ascii ? char_baseaddr_lut_65 : _GEN_1416; // @[CharOutput.scala 118:{17,17}]
  wire [12:0] char_baseaddr_lut_66 = {{1'd0}, _char_baseaddr_lut_T_66}; // @[CharOutput.scala 110:{34,34}]
  wire [12:0] _GEN_1418 = 8'h42 == current_ascii ? char_baseaddr_lut_66 : _GEN_1417; // @[CharOutput.scala 118:{17,17}]
  wire [12:0] char_baseaddr_lut_67 = {{1'd0}, _char_baseaddr_lut_T_67}; // @[CharOutput.scala 110:{34,34}]
  wire [12:0] _GEN_1419 = 8'h43 == current_ascii ? char_baseaddr_lut_67 : _GEN_1418; // @[CharOutput.scala 118:{17,17}]
  wire [12:0] char_baseaddr_lut_68 = {{1'd0}, _char_baseaddr_lut_T_68}; // @[CharOutput.scala 110:{34,34}]
  wire [12:0] _GEN_1420 = 8'h44 == current_ascii ? char_baseaddr_lut_68 : _GEN_1419; // @[CharOutput.scala 118:{17,17}]
  wire [12:0] char_baseaddr_lut_69 = {{1'd0}, _char_baseaddr_lut_T_69}; // @[CharOutput.scala 110:{34,34}]
  wire [12:0] _GEN_1421 = 8'h45 == current_ascii ? char_baseaddr_lut_69 : _GEN_1420; // @[CharOutput.scala 118:{17,17}]
  wire [12:0] char_baseaddr_lut_70 = {{1'd0}, _char_baseaddr_lut_T_70}; // @[CharOutput.scala 110:{34,34}]
  wire [12:0] _GEN_1422 = 8'h46 == current_ascii ? char_baseaddr_lut_70 : _GEN_1421; // @[CharOutput.scala 118:{17,17}]
  wire [12:0] char_baseaddr_lut_71 = {{1'd0}, _char_baseaddr_lut_T_71}; // @[CharOutput.scala 110:{34,34}]
  wire [12:0] _GEN_1423 = 8'h47 == current_ascii ? char_baseaddr_lut_71 : _GEN_1422; // @[CharOutput.scala 118:{17,17}]
  wire [12:0] char_baseaddr_lut_72 = {{1'd0}, _char_baseaddr_lut_T_72}; // @[CharOutput.scala 110:{34,34}]
  wire [12:0] _GEN_1424 = 8'h48 == current_ascii ? char_baseaddr_lut_72 : _GEN_1423; // @[CharOutput.scala 118:{17,17}]
  wire [12:0] char_baseaddr_lut_73 = {{1'd0}, _char_baseaddr_lut_T_73}; // @[CharOutput.scala 110:{34,34}]
  wire [12:0] _GEN_1425 = 8'h49 == current_ascii ? char_baseaddr_lut_73 : _GEN_1424; // @[CharOutput.scala 118:{17,17}]
  wire [12:0] char_baseaddr_lut_74 = {{1'd0}, _char_baseaddr_lut_T_74}; // @[CharOutput.scala 110:{34,34}]
  wire [12:0] _GEN_1426 = 8'h4a == current_ascii ? char_baseaddr_lut_74 : _GEN_1425; // @[CharOutput.scala 118:{17,17}]
  wire [12:0] char_baseaddr_lut_75 = {{1'd0}, _char_baseaddr_lut_T_75}; // @[CharOutput.scala 110:{34,34}]
  wire [12:0] _GEN_1427 = 8'h4b == current_ascii ? char_baseaddr_lut_75 : _GEN_1426; // @[CharOutput.scala 118:{17,17}]
  wire [12:0] char_baseaddr_lut_76 = {{1'd0}, _char_baseaddr_lut_T_76}; // @[CharOutput.scala 110:{34,34}]
  wire [12:0] _GEN_1428 = 8'h4c == current_ascii ? char_baseaddr_lut_76 : _GEN_1427; // @[CharOutput.scala 118:{17,17}]
  wire [12:0] char_baseaddr_lut_77 = {{1'd0}, _char_baseaddr_lut_T_77}; // @[CharOutput.scala 110:{34,34}]
  wire [12:0] _GEN_1429 = 8'h4d == current_ascii ? char_baseaddr_lut_77 : _GEN_1428; // @[CharOutput.scala 118:{17,17}]
  wire [12:0] char_baseaddr_lut_78 = {{1'd0}, _char_baseaddr_lut_T_78}; // @[CharOutput.scala 110:{34,34}]
  wire [12:0] _GEN_1430 = 8'h4e == current_ascii ? char_baseaddr_lut_78 : _GEN_1429; // @[CharOutput.scala 118:{17,17}]
  wire [12:0] char_baseaddr_lut_79 = {{1'd0}, _char_baseaddr_lut_T_79}; // @[CharOutput.scala 110:{34,34}]
  wire [12:0] _GEN_1431 = 8'h4f == current_ascii ? char_baseaddr_lut_79 : _GEN_1430; // @[CharOutput.scala 118:{17,17}]
  wire [12:0] char_baseaddr_lut_80 = {{1'd0}, _char_baseaddr_lut_T_80}; // @[CharOutput.scala 110:{34,34}]
  wire [12:0] _GEN_1432 = 8'h50 == current_ascii ? char_baseaddr_lut_80 : _GEN_1431; // @[CharOutput.scala 118:{17,17}]
  wire [12:0] char_baseaddr_lut_81 = {{1'd0}, _char_baseaddr_lut_T_81}; // @[CharOutput.scala 110:{34,34}]
  wire [12:0] _GEN_1433 = 8'h51 == current_ascii ? char_baseaddr_lut_81 : _GEN_1432; // @[CharOutput.scala 118:{17,17}]
  wire [12:0] char_baseaddr_lut_82 = {{1'd0}, _char_baseaddr_lut_T_82}; // @[CharOutput.scala 110:{34,34}]
  wire [12:0] _GEN_1434 = 8'h52 == current_ascii ? char_baseaddr_lut_82 : _GEN_1433; // @[CharOutput.scala 118:{17,17}]
  wire [12:0] char_baseaddr_lut_83 = {{1'd0}, _char_baseaddr_lut_T_83}; // @[CharOutput.scala 110:{34,34}]
  wire [12:0] _GEN_1435 = 8'h53 == current_ascii ? char_baseaddr_lut_83 : _GEN_1434; // @[CharOutput.scala 118:{17,17}]
  wire [12:0] char_baseaddr_lut_84 = {{1'd0}, _char_baseaddr_lut_T_84}; // @[CharOutput.scala 110:{34,34}]
  wire [12:0] _GEN_1436 = 8'h54 == current_ascii ? char_baseaddr_lut_84 : _GEN_1435; // @[CharOutput.scala 118:{17,17}]
  wire [12:0] char_baseaddr_lut_85 = {{1'd0}, _char_baseaddr_lut_T_85}; // @[CharOutput.scala 110:{34,34}]
  wire [12:0] _GEN_1437 = 8'h55 == current_ascii ? char_baseaddr_lut_85 : _GEN_1436; // @[CharOutput.scala 118:{17,17}]
  wire [12:0] char_baseaddr_lut_86 = {{1'd0}, _char_baseaddr_lut_T_86}; // @[CharOutput.scala 110:{34,34}]
  wire [12:0] _GEN_1438 = 8'h56 == current_ascii ? char_baseaddr_lut_86 : _GEN_1437; // @[CharOutput.scala 118:{17,17}]
  wire [12:0] char_baseaddr_lut_87 = {{1'd0}, _char_baseaddr_lut_T_87}; // @[CharOutput.scala 110:{34,34}]
  wire [12:0] _GEN_1439 = 8'h57 == current_ascii ? char_baseaddr_lut_87 : _GEN_1438; // @[CharOutput.scala 118:{17,17}]
  wire [12:0] char_baseaddr_lut_88 = {{1'd0}, _char_baseaddr_lut_T_88}; // @[CharOutput.scala 110:{34,34}]
  wire [12:0] _GEN_1440 = 8'h58 == current_ascii ? char_baseaddr_lut_88 : _GEN_1439; // @[CharOutput.scala 118:{17,17}]
  wire [12:0] char_baseaddr_lut_89 = {{1'd0}, _char_baseaddr_lut_T_89}; // @[CharOutput.scala 110:{34,34}]
  wire [12:0] _GEN_1441 = 8'h59 == current_ascii ? char_baseaddr_lut_89 : _GEN_1440; // @[CharOutput.scala 118:{17,17}]
  wire [12:0] char_baseaddr_lut_90 = {{1'd0}, _char_baseaddr_lut_T_90}; // @[CharOutput.scala 110:{34,34}]
  wire [12:0] _GEN_1442 = 8'h5a == current_ascii ? char_baseaddr_lut_90 : _GEN_1441; // @[CharOutput.scala 118:{17,17}]
  wire [12:0] char_baseaddr_lut_91 = {{1'd0}, _char_baseaddr_lut_T_91}; // @[CharOutput.scala 110:{34,34}]
  wire [12:0] _GEN_1443 = 8'h5b == current_ascii ? char_baseaddr_lut_91 : _GEN_1442; // @[CharOutput.scala 118:{17,17}]
  wire [12:0] char_baseaddr_lut_92 = {{1'd0}, _char_baseaddr_lut_T_92}; // @[CharOutput.scala 110:{34,34}]
  wire [12:0] _GEN_1444 = 8'h5c == current_ascii ? char_baseaddr_lut_92 : _GEN_1443; // @[CharOutput.scala 118:{17,17}]
  wire [12:0] char_baseaddr_lut_93 = {{1'd0}, _char_baseaddr_lut_T_93}; // @[CharOutput.scala 110:{34,34}]
  wire [12:0] _GEN_1445 = 8'h5d == current_ascii ? char_baseaddr_lut_93 : _GEN_1444; // @[CharOutput.scala 118:{17,17}]
  wire [12:0] char_baseaddr_lut_94 = {{1'd0}, _char_baseaddr_lut_T_94}; // @[CharOutput.scala 110:{34,34}]
  wire [12:0] _GEN_1446 = 8'h5e == current_ascii ? char_baseaddr_lut_94 : _GEN_1445; // @[CharOutput.scala 118:{17,17}]
  wire [12:0] char_baseaddr_lut_95 = {{1'd0}, _char_baseaddr_lut_T_95}; // @[CharOutput.scala 110:{34,34}]
  wire [12:0] _GEN_1447 = 8'h5f == current_ascii ? char_baseaddr_lut_95 : _GEN_1446; // @[CharOutput.scala 118:{17,17}]
  wire [12:0] char_baseaddr_lut_96 = {{1'd0}, _char_baseaddr_lut_T_96}; // @[CharOutput.scala 110:{34,34}]
  wire [12:0] _GEN_1448 = 8'h60 == current_ascii ? char_baseaddr_lut_96 : _GEN_1447; // @[CharOutput.scala 118:{17,17}]
  wire [12:0] char_baseaddr_lut_97 = {{1'd0}, _char_baseaddr_lut_T_97}; // @[CharOutput.scala 110:{34,34}]
  wire [12:0] _GEN_1449 = 8'h61 == current_ascii ? char_baseaddr_lut_97 : _GEN_1448; // @[CharOutput.scala 118:{17,17}]
  wire [12:0] char_baseaddr_lut_98 = {{1'd0}, _char_baseaddr_lut_T_98}; // @[CharOutput.scala 110:{34,34}]
  wire [12:0] _GEN_1450 = 8'h62 == current_ascii ? char_baseaddr_lut_98 : _GEN_1449; // @[CharOutput.scala 118:{17,17}]
  wire [12:0] char_baseaddr_lut_99 = {{1'd0}, _char_baseaddr_lut_T_99}; // @[CharOutput.scala 110:{34,34}]
  wire [12:0] _GEN_1451 = 8'h63 == current_ascii ? char_baseaddr_lut_99 : _GEN_1450; // @[CharOutput.scala 118:{17,17}]
  wire [12:0] char_baseaddr_lut_100 = {{1'd0}, _char_baseaddr_lut_T_100}; // @[CharOutput.scala 110:{34,34}]
  wire [12:0] _GEN_1452 = 8'h64 == current_ascii ? char_baseaddr_lut_100 : _GEN_1451; // @[CharOutput.scala 118:{17,17}]
  wire [12:0] char_baseaddr_lut_101 = {{1'd0}, _char_baseaddr_lut_T_101}; // @[CharOutput.scala 110:{34,34}]
  wire [12:0] _GEN_1453 = 8'h65 == current_ascii ? char_baseaddr_lut_101 : _GEN_1452; // @[CharOutput.scala 118:{17,17}]
  wire [12:0] char_baseaddr_lut_102 = {{1'd0}, _char_baseaddr_lut_T_102}; // @[CharOutput.scala 110:{34,34}]
  wire [12:0] _GEN_1454 = 8'h66 == current_ascii ? char_baseaddr_lut_102 : _GEN_1453; // @[CharOutput.scala 118:{17,17}]
  wire [12:0] char_baseaddr_lut_103 = {{1'd0}, _char_baseaddr_lut_T_103}; // @[CharOutput.scala 110:{34,34}]
  wire [12:0] _GEN_1455 = 8'h67 == current_ascii ? char_baseaddr_lut_103 : _GEN_1454; // @[CharOutput.scala 118:{17,17}]
  wire [12:0] char_baseaddr_lut_104 = {{1'd0}, _char_baseaddr_lut_T_104}; // @[CharOutput.scala 110:{34,34}]
  wire [12:0] _GEN_1456 = 8'h68 == current_ascii ? char_baseaddr_lut_104 : _GEN_1455; // @[CharOutput.scala 118:{17,17}]
  wire [12:0] char_baseaddr_lut_105 = {{1'd0}, _char_baseaddr_lut_T_105}; // @[CharOutput.scala 110:{34,34}]
  wire [12:0] _GEN_1457 = 8'h69 == current_ascii ? char_baseaddr_lut_105 : _GEN_1456; // @[CharOutput.scala 118:{17,17}]
  wire [12:0] char_baseaddr_lut_106 = {{1'd0}, _char_baseaddr_lut_T_106}; // @[CharOutput.scala 110:{34,34}]
  wire [12:0] _GEN_1458 = 8'h6a == current_ascii ? char_baseaddr_lut_106 : _GEN_1457; // @[CharOutput.scala 118:{17,17}]
  wire [12:0] char_baseaddr_lut_107 = {{1'd0}, _char_baseaddr_lut_T_107}; // @[CharOutput.scala 110:{34,34}]
  wire [12:0] _GEN_1459 = 8'h6b == current_ascii ? char_baseaddr_lut_107 : _GEN_1458; // @[CharOutput.scala 118:{17,17}]
  wire [12:0] char_baseaddr_lut_108 = {{1'd0}, _char_baseaddr_lut_T_108}; // @[CharOutput.scala 110:{34,34}]
  wire [12:0] _GEN_1460 = 8'h6c == current_ascii ? char_baseaddr_lut_108 : _GEN_1459; // @[CharOutput.scala 118:{17,17}]
  wire [12:0] char_baseaddr_lut_109 = {{1'd0}, _char_baseaddr_lut_T_109}; // @[CharOutput.scala 110:{34,34}]
  wire [12:0] _GEN_1461 = 8'h6d == current_ascii ? char_baseaddr_lut_109 : _GEN_1460; // @[CharOutput.scala 118:{17,17}]
  wire [12:0] char_baseaddr_lut_110 = {{1'd0}, _char_baseaddr_lut_T_110}; // @[CharOutput.scala 110:{34,34}]
  wire [12:0] _GEN_1462 = 8'h6e == current_ascii ? char_baseaddr_lut_110 : _GEN_1461; // @[CharOutput.scala 118:{17,17}]
  wire [12:0] char_baseaddr_lut_111 = {{1'd0}, _char_baseaddr_lut_T_111}; // @[CharOutput.scala 110:{34,34}]
  wire [12:0] _GEN_1463 = 8'h6f == current_ascii ? char_baseaddr_lut_111 : _GEN_1462; // @[CharOutput.scala 118:{17,17}]
  wire [12:0] char_baseaddr_lut_112 = {{1'd0}, _char_baseaddr_lut_T_112}; // @[CharOutput.scala 110:{34,34}]
  wire [12:0] _GEN_1464 = 8'h70 == current_ascii ? char_baseaddr_lut_112 : _GEN_1463; // @[CharOutput.scala 118:{17,17}]
  wire [12:0] char_baseaddr_lut_113 = {{1'd0}, _char_baseaddr_lut_T_113}; // @[CharOutput.scala 110:{34,34}]
  wire [12:0] _GEN_1465 = 8'h71 == current_ascii ? char_baseaddr_lut_113 : _GEN_1464; // @[CharOutput.scala 118:{17,17}]
  wire [12:0] char_baseaddr_lut_114 = {{1'd0}, _char_baseaddr_lut_T_114}; // @[CharOutput.scala 110:{34,34}]
  wire [12:0] _GEN_1466 = 8'h72 == current_ascii ? char_baseaddr_lut_114 : _GEN_1465; // @[CharOutput.scala 118:{17,17}]
  wire [12:0] char_baseaddr_lut_115 = {{1'd0}, _char_baseaddr_lut_T_115}; // @[CharOutput.scala 110:{34,34}]
  wire [12:0] _GEN_1467 = 8'h73 == current_ascii ? char_baseaddr_lut_115 : _GEN_1466; // @[CharOutput.scala 118:{17,17}]
  wire [12:0] char_baseaddr_lut_116 = {{1'd0}, _char_baseaddr_lut_T_116}; // @[CharOutput.scala 110:{34,34}]
  wire [12:0] _GEN_1468 = 8'h74 == current_ascii ? char_baseaddr_lut_116 : _GEN_1467; // @[CharOutput.scala 118:{17,17}]
  wire [12:0] char_baseaddr_lut_117 = {{1'd0}, _char_baseaddr_lut_T_117}; // @[CharOutput.scala 110:{34,34}]
  wire [12:0] _GEN_1469 = 8'h75 == current_ascii ? char_baseaddr_lut_117 : _GEN_1468; // @[CharOutput.scala 118:{17,17}]
  wire [12:0] char_baseaddr_lut_118 = {{1'd0}, _char_baseaddr_lut_T_118}; // @[CharOutput.scala 110:{34,34}]
  wire [12:0] _GEN_1470 = 8'h76 == current_ascii ? char_baseaddr_lut_118 : _GEN_1469; // @[CharOutput.scala 118:{17,17}]
  wire [12:0] char_baseaddr_lut_119 = {{1'd0}, _char_baseaddr_lut_T_119}; // @[CharOutput.scala 110:{34,34}]
  wire [12:0] _GEN_1471 = 8'h77 == current_ascii ? char_baseaddr_lut_119 : _GEN_1470; // @[CharOutput.scala 118:{17,17}]
  wire [12:0] char_baseaddr_lut_120 = {{1'd0}, _char_baseaddr_lut_T_120}; // @[CharOutput.scala 110:{34,34}]
  wire [12:0] _GEN_1472 = 8'h78 == current_ascii ? char_baseaddr_lut_120 : _GEN_1471; // @[CharOutput.scala 118:{17,17}]
  wire [12:0] char_baseaddr_lut_121 = {{1'd0}, _char_baseaddr_lut_T_121}; // @[CharOutput.scala 110:{34,34}]
  wire [12:0] _GEN_1473 = 8'h79 == current_ascii ? char_baseaddr_lut_121 : _GEN_1472; // @[CharOutput.scala 118:{17,17}]
  wire [12:0] char_baseaddr_lut_122 = {{1'd0}, _char_baseaddr_lut_T_122}; // @[CharOutput.scala 110:{34,34}]
  wire [12:0] _GEN_1474 = 8'h7a == current_ascii ? char_baseaddr_lut_122 : _GEN_1473; // @[CharOutput.scala 118:{17,17}]
  wire [12:0] char_baseaddr_lut_123 = {{1'd0}, _char_baseaddr_lut_T_123}; // @[CharOutput.scala 110:{34,34}]
  wire [12:0] _GEN_1475 = 8'h7b == current_ascii ? char_baseaddr_lut_123 : _GEN_1474; // @[CharOutput.scala 118:{17,17}]
  wire [12:0] char_baseaddr_lut_124 = {{1'd0}, _char_baseaddr_lut_T_124}; // @[CharOutput.scala 110:{34,34}]
  wire [12:0] _GEN_1476 = 8'h7c == current_ascii ? char_baseaddr_lut_124 : _GEN_1475; // @[CharOutput.scala 118:{17,17}]
  wire [12:0] char_baseaddr_lut_125 = {{1'd0}, _char_baseaddr_lut_T_125}; // @[CharOutput.scala 110:{34,34}]
  wire [12:0] _GEN_1477 = 8'h7d == current_ascii ? char_baseaddr_lut_125 : _GEN_1476; // @[CharOutput.scala 118:{17,17}]
  wire [12:0] char_baseaddr_lut_126 = {{1'd0}, _char_baseaddr_lut_T_126}; // @[CharOutput.scala 110:{34,34}]
  wire [12:0] _GEN_1478 = 8'h7e == current_ascii ? char_baseaddr_lut_126 : _GEN_1477; // @[CharOutput.scala 118:{17,17}]
  wire [12:0] char_baseaddr_lut_127 = {{1'd0}, _char_baseaddr_lut_T_127}; // @[CharOutput.scala 110:{34,34}]
  wire [12:0] _GEN_1479 = 8'h7f == current_ascii ? char_baseaddr_lut_127 : _GEN_1478; // @[CharOutput.scala 118:{17,17}]
  wire [12:0] _GEN_1480 = 8'h80 == current_ascii ? char_baseaddr_lut_128 : _GEN_1479; // @[CharOutput.scala 118:{17,17}]
  wire [12:0] _GEN_1481 = 8'h81 == current_ascii ? char_baseaddr_lut_129 : _GEN_1480; // @[CharOutput.scala 118:{17,17}]
  wire [12:0] _GEN_1482 = 8'h82 == current_ascii ? char_baseaddr_lut_130 : _GEN_1481; // @[CharOutput.scala 118:{17,17}]
  wire [12:0] _GEN_1483 = 8'h83 == current_ascii ? char_baseaddr_lut_131 : _GEN_1482; // @[CharOutput.scala 118:{17,17}]
  wire [12:0] _GEN_1484 = 8'h84 == current_ascii ? char_baseaddr_lut_132 : _GEN_1483; // @[CharOutput.scala 118:{17,17}]
  wire [12:0] _GEN_1485 = 8'h85 == current_ascii ? char_baseaddr_lut_133 : _GEN_1484; // @[CharOutput.scala 118:{17,17}]
  wire [12:0] _GEN_1486 = 8'h86 == current_ascii ? char_baseaddr_lut_134 : _GEN_1485; // @[CharOutput.scala 118:{17,17}]
  wire [12:0] _GEN_1487 = 8'h87 == current_ascii ? char_baseaddr_lut_135 : _GEN_1486; // @[CharOutput.scala 118:{17,17}]
  wire [12:0] _GEN_1488 = 8'h88 == current_ascii ? char_baseaddr_lut_136 : _GEN_1487; // @[CharOutput.scala 118:{17,17}]
  wire [12:0] _GEN_1489 = 8'h89 == current_ascii ? char_baseaddr_lut_137 : _GEN_1488; // @[CharOutput.scala 118:{17,17}]
  wire [12:0] _GEN_1490 = 8'h8a == current_ascii ? char_baseaddr_lut_138 : _GEN_1489; // @[CharOutput.scala 118:{17,17}]
  wire [12:0] _GEN_1491 = 8'h8b == current_ascii ? char_baseaddr_lut_139 : _GEN_1490; // @[CharOutput.scala 118:{17,17}]
  wire [12:0] _GEN_1492 = 8'h8c == current_ascii ? char_baseaddr_lut_140 : _GEN_1491; // @[CharOutput.scala 118:{17,17}]
  wire [12:0] _GEN_1493 = 8'h8d == current_ascii ? char_baseaddr_lut_141 : _GEN_1492; // @[CharOutput.scala 118:{17,17}]
  wire [12:0] _GEN_1494 = 8'h8e == current_ascii ? char_baseaddr_lut_142 : _GEN_1493; // @[CharOutput.scala 118:{17,17}]
  wire [12:0] _GEN_1495 = 8'h8f == current_ascii ? char_baseaddr_lut_143 : _GEN_1494; // @[CharOutput.scala 118:{17,17}]
  wire [12:0] _GEN_1496 = 8'h90 == current_ascii ? char_baseaddr_lut_144 : _GEN_1495; // @[CharOutput.scala 118:{17,17}]
  wire [12:0] _GEN_1497 = 8'h91 == current_ascii ? char_baseaddr_lut_145 : _GEN_1496; // @[CharOutput.scala 118:{17,17}]
  wire [12:0] _GEN_1498 = 8'h92 == current_ascii ? char_baseaddr_lut_146 : _GEN_1497; // @[CharOutput.scala 118:{17,17}]
  wire [12:0] _GEN_1499 = 8'h93 == current_ascii ? char_baseaddr_lut_147 : _GEN_1498; // @[CharOutput.scala 118:{17,17}]
  wire [12:0] _GEN_1500 = 8'h94 == current_ascii ? char_baseaddr_lut_148 : _GEN_1499; // @[CharOutput.scala 118:{17,17}]
  wire [12:0] _GEN_1501 = 8'h95 == current_ascii ? char_baseaddr_lut_149 : _GEN_1500; // @[CharOutput.scala 118:{17,17}]
  wire [12:0] _GEN_1502 = 8'h96 == current_ascii ? char_baseaddr_lut_150 : _GEN_1501; // @[CharOutput.scala 118:{17,17}]
  wire [12:0] _GEN_1503 = 8'h97 == current_ascii ? char_baseaddr_lut_151 : _GEN_1502; // @[CharOutput.scala 118:{17,17}]
  wire [12:0] _GEN_1504 = 8'h98 == current_ascii ? char_baseaddr_lut_152 : _GEN_1503; // @[CharOutput.scala 118:{17,17}]
  wire [12:0] _GEN_1505 = 8'h99 == current_ascii ? char_baseaddr_lut_153 : _GEN_1504; // @[CharOutput.scala 118:{17,17}]
  wire [12:0] _GEN_1506 = 8'h9a == current_ascii ? char_baseaddr_lut_154 : _GEN_1505; // @[CharOutput.scala 118:{17,17}]
  wire [12:0] _GEN_1507 = 8'h9b == current_ascii ? char_baseaddr_lut_155 : _GEN_1506; // @[CharOutput.scala 118:{17,17}]
  wire [12:0] _GEN_1508 = 8'h9c == current_ascii ? char_baseaddr_lut_156 : _GEN_1507; // @[CharOutput.scala 118:{17,17}]
  wire [12:0] _GEN_1509 = 8'h9d == current_ascii ? char_baseaddr_lut_157 : _GEN_1508; // @[CharOutput.scala 118:{17,17}]
  wire [12:0] _GEN_1510 = 8'h9e == current_ascii ? char_baseaddr_lut_158 : _GEN_1509; // @[CharOutput.scala 118:{17,17}]
  wire [12:0] _GEN_1511 = 8'h9f == current_ascii ? char_baseaddr_lut_159 : _GEN_1510; // @[CharOutput.scala 118:{17,17}]
  wire [12:0] _GEN_1512 = 8'ha0 == current_ascii ? char_baseaddr_lut_160 : _GEN_1511; // @[CharOutput.scala 118:{17,17}]
  wire [12:0] _GEN_1513 = 8'ha1 == current_ascii ? char_baseaddr_lut_161 : _GEN_1512; // @[CharOutput.scala 118:{17,17}]
  wire [12:0] _GEN_1514 = 8'ha2 == current_ascii ? char_baseaddr_lut_162 : _GEN_1513; // @[CharOutput.scala 118:{17,17}]
  wire [12:0] _GEN_1515 = 8'ha3 == current_ascii ? char_baseaddr_lut_163 : _GEN_1514; // @[CharOutput.scala 118:{17,17}]
  wire [12:0] _GEN_1516 = 8'ha4 == current_ascii ? char_baseaddr_lut_164 : _GEN_1515; // @[CharOutput.scala 118:{17,17}]
  wire [12:0] _GEN_1517 = 8'ha5 == current_ascii ? char_baseaddr_lut_165 : _GEN_1516; // @[CharOutput.scala 118:{17,17}]
  wire [12:0] _GEN_1518 = 8'ha6 == current_ascii ? char_baseaddr_lut_166 : _GEN_1517; // @[CharOutput.scala 118:{17,17}]
  wire [12:0] _GEN_1519 = 8'ha7 == current_ascii ? char_baseaddr_lut_167 : _GEN_1518; // @[CharOutput.scala 118:{17,17}]
  wire [12:0] _GEN_1520 = 8'ha8 == current_ascii ? char_baseaddr_lut_168 : _GEN_1519; // @[CharOutput.scala 118:{17,17}]
  wire [12:0] _GEN_1521 = 8'ha9 == current_ascii ? char_baseaddr_lut_169 : _GEN_1520; // @[CharOutput.scala 118:{17,17}]
  wire [12:0] _GEN_1522 = 8'haa == current_ascii ? char_baseaddr_lut_170 : _GEN_1521; // @[CharOutput.scala 118:{17,17}]
  wire [12:0] _GEN_1523 = 8'hab == current_ascii ? char_baseaddr_lut_171 : _GEN_1522; // @[CharOutput.scala 118:{17,17}]
  wire [12:0] _GEN_1524 = 8'hac == current_ascii ? char_baseaddr_lut_172 : _GEN_1523; // @[CharOutput.scala 118:{17,17}]
  wire [12:0] _GEN_1525 = 8'had == current_ascii ? char_baseaddr_lut_173 : _GEN_1524; // @[CharOutput.scala 118:{17,17}]
  wire [12:0] _GEN_1526 = 8'hae == current_ascii ? char_baseaddr_lut_174 : _GEN_1525; // @[CharOutput.scala 118:{17,17}]
  wire [12:0] _GEN_1527 = 8'haf == current_ascii ? char_baseaddr_lut_175 : _GEN_1526; // @[CharOutput.scala 118:{17,17}]
  wire [12:0] _GEN_1528 = 8'hb0 == current_ascii ? char_baseaddr_lut_176 : _GEN_1527; // @[CharOutput.scala 118:{17,17}]
  wire [12:0] _GEN_1529 = 8'hb1 == current_ascii ? char_baseaddr_lut_177 : _GEN_1528; // @[CharOutput.scala 118:{17,17}]
  wire [12:0] _GEN_1530 = 8'hb2 == current_ascii ? char_baseaddr_lut_178 : _GEN_1529; // @[CharOutput.scala 118:{17,17}]
  wire [12:0] _GEN_1531 = 8'hb3 == current_ascii ? char_baseaddr_lut_179 : _GEN_1530; // @[CharOutput.scala 118:{17,17}]
  wire [12:0] _GEN_1532 = 8'hb4 == current_ascii ? char_baseaddr_lut_180 : _GEN_1531; // @[CharOutput.scala 118:{17,17}]
  wire [12:0] _GEN_1533 = 8'hb5 == current_ascii ? char_baseaddr_lut_181 : _GEN_1532; // @[CharOutput.scala 118:{17,17}]
  wire [12:0] _GEN_1534 = 8'hb6 == current_ascii ? char_baseaddr_lut_182 : _GEN_1533; // @[CharOutput.scala 118:{17,17}]
  wire [12:0] _GEN_1535 = 8'hb7 == current_ascii ? char_baseaddr_lut_183 : _GEN_1534; // @[CharOutput.scala 118:{17,17}]
  wire [12:0] _GEN_1536 = 8'hb8 == current_ascii ? char_baseaddr_lut_184 : _GEN_1535; // @[CharOutput.scala 118:{17,17}]
  wire [12:0] _GEN_1537 = 8'hb9 == current_ascii ? char_baseaddr_lut_185 : _GEN_1536; // @[CharOutput.scala 118:{17,17}]
  wire [12:0] _GEN_1538 = 8'hba == current_ascii ? char_baseaddr_lut_186 : _GEN_1537; // @[CharOutput.scala 118:{17,17}]
  wire [12:0] _GEN_1539 = 8'hbb == current_ascii ? char_baseaddr_lut_187 : _GEN_1538; // @[CharOutput.scala 118:{17,17}]
  wire [12:0] _GEN_1540 = 8'hbc == current_ascii ? char_baseaddr_lut_188 : _GEN_1539; // @[CharOutput.scala 118:{17,17}]
  wire [12:0] _GEN_1541 = 8'hbd == current_ascii ? char_baseaddr_lut_189 : _GEN_1540; // @[CharOutput.scala 118:{17,17}]
  wire [12:0] _GEN_1542 = 8'hbe == current_ascii ? char_baseaddr_lut_190 : _GEN_1541; // @[CharOutput.scala 118:{17,17}]
  wire [12:0] _GEN_1543 = 8'hbf == current_ascii ? char_baseaddr_lut_191 : _GEN_1542; // @[CharOutput.scala 118:{17,17}]
  wire [12:0] _GEN_1544 = 8'hc0 == current_ascii ? char_baseaddr_lut_192 : _GEN_1543; // @[CharOutput.scala 118:{17,17}]
  wire [12:0] _GEN_1545 = 8'hc1 == current_ascii ? char_baseaddr_lut_193 : _GEN_1544; // @[CharOutput.scala 118:{17,17}]
  wire [12:0] _GEN_1546 = 8'hc2 == current_ascii ? char_baseaddr_lut_194 : _GEN_1545; // @[CharOutput.scala 118:{17,17}]
  wire [12:0] _GEN_1547 = 8'hc3 == current_ascii ? char_baseaddr_lut_195 : _GEN_1546; // @[CharOutput.scala 118:{17,17}]
  wire [12:0] _GEN_1548 = 8'hc4 == current_ascii ? char_baseaddr_lut_196 : _GEN_1547; // @[CharOutput.scala 118:{17,17}]
  wire [12:0] _GEN_1549 = 8'hc5 == current_ascii ? char_baseaddr_lut_197 : _GEN_1548; // @[CharOutput.scala 118:{17,17}]
  wire [12:0] _GEN_1550 = 8'hc6 == current_ascii ? char_baseaddr_lut_198 : _GEN_1549; // @[CharOutput.scala 118:{17,17}]
  wire [12:0] _GEN_1551 = 8'hc7 == current_ascii ? char_baseaddr_lut_199 : _GEN_1550; // @[CharOutput.scala 118:{17,17}]
  wire [12:0] _GEN_1552 = 8'hc8 == current_ascii ? char_baseaddr_lut_200 : _GEN_1551; // @[CharOutput.scala 118:{17,17}]
  wire [12:0] _GEN_1553 = 8'hc9 == current_ascii ? char_baseaddr_lut_201 : _GEN_1552; // @[CharOutput.scala 118:{17,17}]
  wire [12:0] _GEN_1554 = 8'hca == current_ascii ? char_baseaddr_lut_202 : _GEN_1553; // @[CharOutput.scala 118:{17,17}]
  wire [12:0] _GEN_1555 = 8'hcb == current_ascii ? char_baseaddr_lut_203 : _GEN_1554; // @[CharOutput.scala 118:{17,17}]
  wire [12:0] _GEN_1556 = 8'hcc == current_ascii ? char_baseaddr_lut_204 : _GEN_1555; // @[CharOutput.scala 118:{17,17}]
  wire [12:0] _GEN_1557 = 8'hcd == current_ascii ? char_baseaddr_lut_205 : _GEN_1556; // @[CharOutput.scala 118:{17,17}]
  wire [12:0] _GEN_1558 = 8'hce == current_ascii ? char_baseaddr_lut_206 : _GEN_1557; // @[CharOutput.scala 118:{17,17}]
  wire [12:0] _GEN_1559 = 8'hcf == current_ascii ? char_baseaddr_lut_207 : _GEN_1558; // @[CharOutput.scala 118:{17,17}]
  wire [12:0] _GEN_1560 = 8'hd0 == current_ascii ? char_baseaddr_lut_208 : _GEN_1559; // @[CharOutput.scala 118:{17,17}]
  wire [12:0] _GEN_1561 = 8'hd1 == current_ascii ? char_baseaddr_lut_209 : _GEN_1560; // @[CharOutput.scala 118:{17,17}]
  wire [12:0] _GEN_1562 = 8'hd2 == current_ascii ? char_baseaddr_lut_210 : _GEN_1561; // @[CharOutput.scala 118:{17,17}]
  wire [12:0] _GEN_1563 = 8'hd3 == current_ascii ? char_baseaddr_lut_211 : _GEN_1562; // @[CharOutput.scala 118:{17,17}]
  wire [12:0] _GEN_1564 = 8'hd4 == current_ascii ? char_baseaddr_lut_212 : _GEN_1563; // @[CharOutput.scala 118:{17,17}]
  wire [12:0] _GEN_1565 = 8'hd5 == current_ascii ? char_baseaddr_lut_213 : _GEN_1564; // @[CharOutput.scala 118:{17,17}]
  wire [12:0] _GEN_1566 = 8'hd6 == current_ascii ? char_baseaddr_lut_214 : _GEN_1565; // @[CharOutput.scala 118:{17,17}]
  wire [12:0] _GEN_1567 = 8'hd7 == current_ascii ? char_baseaddr_lut_215 : _GEN_1566; // @[CharOutput.scala 118:{17,17}]
  wire [12:0] _GEN_1568 = 8'hd8 == current_ascii ? char_baseaddr_lut_216 : _GEN_1567; // @[CharOutput.scala 118:{17,17}]
  wire [12:0] _GEN_1569 = 8'hd9 == current_ascii ? char_baseaddr_lut_217 : _GEN_1568; // @[CharOutput.scala 118:{17,17}]
  wire [12:0] _GEN_1570 = 8'hda == current_ascii ? char_baseaddr_lut_218 : _GEN_1569; // @[CharOutput.scala 118:{17,17}]
  wire [12:0] _GEN_1571 = 8'hdb == current_ascii ? char_baseaddr_lut_219 : _GEN_1570; // @[CharOutput.scala 118:{17,17}]
  wire [12:0] _GEN_1572 = 8'hdc == current_ascii ? char_baseaddr_lut_220 : _GEN_1571; // @[CharOutput.scala 118:{17,17}]
  wire [12:0] _GEN_1573 = 8'hdd == current_ascii ? char_baseaddr_lut_221 : _GEN_1572; // @[CharOutput.scala 118:{17,17}]
  wire [12:0] _GEN_1574 = 8'hde == current_ascii ? char_baseaddr_lut_222 : _GEN_1573; // @[CharOutput.scala 118:{17,17}]
  wire [12:0] _GEN_1575 = 8'hdf == current_ascii ? char_baseaddr_lut_223 : _GEN_1574; // @[CharOutput.scala 118:{17,17}]
  wire [12:0] _GEN_1576 = 8'he0 == current_ascii ? char_baseaddr_lut_224 : _GEN_1575; // @[CharOutput.scala 118:{17,17}]
  wire [12:0] _GEN_1577 = 8'he1 == current_ascii ? char_baseaddr_lut_225 : _GEN_1576; // @[CharOutput.scala 118:{17,17}]
  wire [12:0] _GEN_1578 = 8'he2 == current_ascii ? char_baseaddr_lut_226 : _GEN_1577; // @[CharOutput.scala 118:{17,17}]
  wire [12:0] _GEN_1579 = 8'he3 == current_ascii ? char_baseaddr_lut_227 : _GEN_1578; // @[CharOutput.scala 118:{17,17}]
  wire [12:0] _GEN_1580 = 8'he4 == current_ascii ? char_baseaddr_lut_228 : _GEN_1579; // @[CharOutput.scala 118:{17,17}]
  wire [12:0] _GEN_1581 = 8'he5 == current_ascii ? char_baseaddr_lut_229 : _GEN_1580; // @[CharOutput.scala 118:{17,17}]
  wire [12:0] _GEN_1582 = 8'he6 == current_ascii ? char_baseaddr_lut_230 : _GEN_1581; // @[CharOutput.scala 118:{17,17}]
  wire [12:0] _GEN_1583 = 8'he7 == current_ascii ? char_baseaddr_lut_231 : _GEN_1582; // @[CharOutput.scala 118:{17,17}]
  wire [12:0] _GEN_1584 = 8'he8 == current_ascii ? char_baseaddr_lut_232 : _GEN_1583; // @[CharOutput.scala 118:{17,17}]
  wire [12:0] _GEN_1585 = 8'he9 == current_ascii ? char_baseaddr_lut_233 : _GEN_1584; // @[CharOutput.scala 118:{17,17}]
  wire [12:0] _GEN_1586 = 8'hea == current_ascii ? char_baseaddr_lut_234 : _GEN_1585; // @[CharOutput.scala 118:{17,17}]
  wire [12:0] _GEN_1587 = 8'heb == current_ascii ? char_baseaddr_lut_235 : _GEN_1586; // @[CharOutput.scala 118:{17,17}]
  wire [12:0] _GEN_1588 = 8'hec == current_ascii ? char_baseaddr_lut_236 : _GEN_1587; // @[CharOutput.scala 118:{17,17}]
  wire [12:0] _GEN_1589 = 8'hed == current_ascii ? char_baseaddr_lut_237 : _GEN_1588; // @[CharOutput.scala 118:{17,17}]
  wire [12:0] _GEN_1590 = 8'hee == current_ascii ? char_baseaddr_lut_238 : _GEN_1589; // @[CharOutput.scala 118:{17,17}]
  wire [12:0] _GEN_1591 = 8'hef == current_ascii ? char_baseaddr_lut_239 : _GEN_1590; // @[CharOutput.scala 118:{17,17}]
  wire [12:0] _GEN_1592 = 8'hf0 == current_ascii ? char_baseaddr_lut_240 : _GEN_1591; // @[CharOutput.scala 118:{17,17}]
  wire [12:0] _GEN_1593 = 8'hf1 == current_ascii ? char_baseaddr_lut_241 : _GEN_1592; // @[CharOutput.scala 118:{17,17}]
  wire [12:0] _GEN_1594 = 8'hf2 == current_ascii ? char_baseaddr_lut_242 : _GEN_1593; // @[CharOutput.scala 118:{17,17}]
  wire [12:0] _GEN_1595 = 8'hf3 == current_ascii ? char_baseaddr_lut_243 : _GEN_1594; // @[CharOutput.scala 118:{17,17}]
  wire [12:0] _GEN_1596 = 8'hf4 == current_ascii ? char_baseaddr_lut_244 : _GEN_1595; // @[CharOutput.scala 118:{17,17}]
  wire [12:0] _GEN_1597 = 8'hf5 == current_ascii ? char_baseaddr_lut_245 : _GEN_1596; // @[CharOutput.scala 118:{17,17}]
  wire [12:0] _GEN_1598 = 8'hf6 == current_ascii ? char_baseaddr_lut_246 : _GEN_1597; // @[CharOutput.scala 118:{17,17}]
  wire [12:0] _GEN_1599 = 8'hf7 == current_ascii ? char_baseaddr_lut_247 : _GEN_1598; // @[CharOutput.scala 118:{17,17}]
  wire [12:0] _GEN_1600 = 8'hf8 == current_ascii ? char_baseaddr_lut_248 : _GEN_1599; // @[CharOutput.scala 118:{17,17}]
  wire [12:0] _GEN_1601 = 8'hf9 == current_ascii ? char_baseaddr_lut_249 : _GEN_1600; // @[CharOutput.scala 118:{17,17}]
  wire [12:0] _GEN_1602 = 8'hfa == current_ascii ? char_baseaddr_lut_250 : _GEN_1601; // @[CharOutput.scala 118:{17,17}]
  wire [12:0] _GEN_1603 = 8'hfb == current_ascii ? char_baseaddr_lut_251 : _GEN_1602; // @[CharOutput.scala 118:{17,17}]
  wire [12:0] _GEN_1604 = 8'hfc == current_ascii ? char_baseaddr_lut_252 : _GEN_1603; // @[CharOutput.scala 118:{17,17}]
  wire [12:0] _GEN_1605 = 8'hfd == current_ascii ? char_baseaddr_lut_253 : _GEN_1604; // @[CharOutput.scala 118:{17,17}]
  wire [12:0] _GEN_1606 = 8'hfe == current_ascii ? char_baseaddr_lut_254 : _GEN_1605; // @[CharOutput.scala 118:{17,17}]
  wire [12:0] char_baseaddr = 8'hff == current_ascii ? char_baseaddr_lut_255 : _GEN_1606; // @[CharOutput.scala 118:{17,17}]
  wire [3:0] char_row_0 = _GEN_305[3:0]; // @[CharOutput.scala 76:25]
  wire [3:0] char_row_1 = _GEN_506[3:0]; // @[CharOutput.scala 76:25]
  wire [3:0] _GEN_1609 = 3'h1 == obj_choose ? char_row_1 : char_row_0; // @[CharOutput.scala 119:{31,31}]
  wire [3:0] char_row_2 = _GEN_707[3:0]; // @[CharOutput.scala 76:25]
  wire [3:0] _GEN_1610 = 3'h2 == obj_choose ? char_row_2 : _GEN_1609; // @[CharOutput.scala 119:{31,31}]
  wire [3:0] char_row_3 = _GEN_908[3:0]; // @[CharOutput.scala 76:25]
  wire [3:0] _GEN_1611 = 3'h3 == obj_choose ? char_row_3 : _GEN_1610; // @[CharOutput.scala 119:{31,31}]
  wire [3:0] char_row_4 = _GEN_1109[3:0]; // @[CharOutput.scala 76:25]
  wire [3:0] _GEN_1612 = 3'h4 == obj_choose ? char_row_4 : _GEN_1611; // @[CharOutput.scala 119:{31,31}]
  wire [12:0] _GEN_1623 = {{9'd0}, _GEN_1612}; // @[CharOutput.scala 119:31]
  wire [12:0] piexl_addr = char_baseaddr + _GEN_1623; // @[CharOutput.scala 119:31]
  wire [3:0] _GEN_1614 = 3'h1 == obj_choose ? char_col_1 : char_col_0; // @[CharOutput.scala 120:{35,35}]
  wire [3:0] _GEN_1615 = 3'h2 == obj_choose ? char_col_2 : _GEN_1614; // @[CharOutput.scala 120:{35,35}]
  wire [3:0] _GEN_1616 = 3'h3 == obj_choose ? char_col_3 : _GEN_1615; // @[CharOutput.scala 120:{35,35}]
  wire [3:0] _GEN_1617 = 3'h4 == obj_choose ? char_col_4 : _GEN_1616; // @[CharOutput.scala 120:{35,35}]
  wire [11:0] _io_pixel_T_2 = dot_txt_io_pixel_MPORT_data >> _GEN_1617; // @[CharOutput.scala 120:35]
  assign dot_txt_io_pixel_MPORT_en = 1'h1;
  assign dot_txt_io_pixel_MPORT_addr = piexl_addr[11:0];
  assign dot_txt_io_pixel_MPORT_data = dot_txt[dot_txt_io_pixel_MPORT_addr]; // @[CharOutput.scala 105:20]
  assign io_pixel = _io_pixel_T_2[0] & _T_11; // @[CharOutput.scala 120:66]
  assign io_char_area_valid_0 = enc[0]; // @[OneHot.scala 82:30]
  assign io_char_area_valid_1 = enc[1]; // @[OneHot.scala 82:30]
  assign io_char_area_valid_2 = enc[2]; // @[OneHot.scala 82:30]
  assign io_char_area_valid_3 = enc[3]; // @[OneHot.scala 82:30]
  assign io_char_area_valid_4 = enc[4]; // @[OneHot.scala 82:30]

initial begin
  $readmemh("C:/Users/Administrator/Desktop/jichuang_code_7_12/font_txt.txt", dot_txt);
end // initial

endmodule
